--------------------------------------------------------------------------------
-- This file is part of the ParaNut project.
-- 
-- Copyright (C) 2013  Michael Seider, Hochschule Augsburg
-- michael.seider@hs-augsburg.de
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
-- Description:
--  Readport module for the MEMU.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library paranut;
use paranut.paranut_config.all;
use paranut.types.all;
use paranut.memu_lib.all;
use paranut.paranut_lib.all;
use paranut.histogram.all;

entity mwriteport is
    port (
             clk    : in std_logic;
             reset  : in std_logic;
             -- With (CPU) port...
             wpi    : in writeport_in_type;
             wpo    : out writeport_out_type;
             -- With cache...
             wpci   : in writeport_cache_in_type;
             wpco   : out writeport_cache_out_type;
             -- With BUSIF...
             wpbifi : in writeport_busif_in_type;
             wpbifo : out writeport_busif_out_type;
             -- Request & grant lines...
             wpai   : in writeport_arbiter_in_type;
             wpao   : out writeport_arbiter_out_type;
             -- Histogram...
             hist_cache_write_hit : out hist_ctrl_type;
             hist_cache_write_miss : out hist_ctrl_type
         );
end mwriteport;

architecture rtl of mwriteport is

-- - All input ports must be held until 'port_ack' is asserted, at least for one cycle.
-- - 'port_ack' is issued for exactly one cycle (no full handshake).
-- - 'port_ack' may be asserted already in the same cycle as the request was issued.
-- - The next request may be issued at earliest one cycle after 'port_ack' was asserted (TBD: allow in the ACK cycle?)
-- - If 'port_direct' is set, nothing happens with the cache (i.e. no invalidation).
--   Hence, 'port_direct' = 0/1 should not be mixed for one address.

    type state_type is (S_WP_INIT, S_WP_DIRECT, S_WP_REQUEST_LINELOCK_ONLY,
    S_WP_READ_TAG, S_WP_HAVE_TAG_REQUEST_BANK, S_WP_READ_BANK,
    S_WP_WRITE_TAG1_AND_BANK, S_WP_WRITE_TAG2_AND_BANK, S_WP_WRITE_TAG1,
    S_WP_WRITE_TAG2, S_WP_WRITE_BANK, S_WP_MISS, S_WP_REQUEST_BUSIF_ONLY,
    S_WP_RECHECK, S_WP_RECHECK_READ_TAG, S_WP_REPLACE, S_WP_REPLACE_WAIT_BUSIF,
    S_WP_SPECIAL_REQUEST_BUSIF_ONLY, S_WP_SPECIAL, S_WP_SPECIAL_WAIT_COMPLETE);

    function combine_data (bsel : TByteSel; word0, word1 : TWord) return TWord
    is
        variable ret : TWord;
    begin
        ret := word1;
        for n in 0 to 3 loop
            if (bsel(3-n) = '0') then
                ret(8*(n+1)-1 downto 8*n) := word0(8*(n+1)-1 downto 8*n);
            end if;
        end loop;
        return (ret);
    end;

    type registers is record
        state : state_type;
        tag : cache_tag_type;
        data : TWord;
        link_adr : TWord;
        link_valid : std_logic;
        -- Histogram...
        hist_miss : std_logic;
    end record;

    signal r, rin : registers;

begin

    comb : process (r, reset, wpi, wpbifi, wpci, wpai)
        variable v : registers;
        -- Output variables
        variable vwpo : writeport_out_type;
        variable vwpbifo : writeport_busif_out_type;
        variable vwpco : writeport_cache_out_type;
        variable vwpao : writeport_arbiter_out_type;
        -- Helper variables
        variable tag : cache_tag_type;
        variable index : std_logic_vector(CFG_MEMU_CACHE_SETS_LD-1 downto 0);
        variable bank : std_logic_vector(CFG_MEMU_CACHE_BANKS_LD-1 downto 0);
        variable data : TWord;
        variable bank_req_rd : std_logic;
        variable bank_gnt : std_logic;
    begin

        v := r;
        -- Defaults for outputs...

        hist_cache_write_hit.start <= '0';
        hist_cache_write_hit.stop <= '0';
        hist_cache_write_hit.abort <= '0';
        hist_cache_write_miss.start <= '0';
        hist_cache_write_miss.stop <= '0';
        hist_cache_write_miss.abort <= '0';

        vwpo.port_ack := '0';
        vwpo.port_wcond_ok := r.link_valid;

        vwpbifo.busif_op := BIO_NOTHING;
        vwpbifo.busif_nolinelock := '1';

        vwpco.tag_rd := '0';
        vwpco.tag_wr := '0';
        vwpco.bank_wr := '0';
        vwpco.tag_out := r.tag;
        --vwpco.bank_data_out := (others => '-'); --TODO
        vwpco.bank_data_out := combine_data(wpi.port_bsel, r.data, wpi.port_data);

        vwpao.req_linelock := '0';
        vwpao.req_tagr := '0';
        vwpao.req_tagw := '0';
        vwpao.req_bank := (others => '0');
        vwpao.req_busif := '0';

        -- Helper variables
        index := wpi.port_adr(INDEX_OF_ADDR_RANGE);
        bank := wpi.port_adr(BANK_OF_ADDR_RANGE);
        bank_req_rd := '0';
        bank_gnt := wpai.gnt_bank(conv_integer(bank));

        -- Update link registers...
        if (wpai.snoop_stb = '1') then
            if (wpai.snoop_adr = r.link_adr) then -- need to invalidate?
                v.link_valid := '0';
            end if;
        end if;

        -- Main "switch"...
        if (reset = '1') then
            v.state := S_WP_INIT;
            v.link_valid := '0';
        else
            case r.state is
                when S_WP_INIT =>
                    if (wpi.port_wr = '1') then
                        if (wpi.port_direct = '1') then
                            -- Direct (uncached) memory access...
                            vwpao.req_busif := '1';
                            vwpbifo.busif_op := BIO_DIRECT_WRITE;
                            if (wpai.gnt_busif = '1' and wpbifi.busif_busy = '0') then
                                v.state := S_WP_DIRECT;
                            end if;
                        else
                            -- Normal (cached) access...
                            if (wpi.port_rlink_wcond = '1' and r.link_valid = '0') then
                                -- This is a "store conditional" (SC), which has failed right away...
                                -- (a failure may still occur later, even if this condition has not yet been fulfilled here)
                                vwpo.port_ack := '1';
                            else
                                -- Normal and (so far) successful SC cache accesses...
                                if (CFG_NUT_HISTOGRAM) then
                                    v.hist_miss := '0';
                                end if;
                                hist_cache_write_hit.start <= '1';
                                hist_cache_write_miss.start <= '1';
                                vwpao.req_linelock := '1';
                                vwpao.req_tagr := '1';
                                if (wpai.gnt_tagr = '1') then
                                    vwpco.tag_rd := '1';
                                    if (wpai.gnt_linelock = '1') then
                                        v.state := S_WP_READ_TAG;
                                    else
                                        v.state := S_WP_REQUEST_LINELOCK_ONLY;
                                    end if;
                                end if;
                            end if;
                        end if;
                    elsif (wpi.port_writeback = '1' or wpi.port_invalidate = '1') then
                        -- Special operation...
                        vwpao.req_busif := '1';
                        vwpao.req_linelock := '1';
                        if (wpai.gnt_linelock = '1' and wpai.gnt_busif = '0') then
                            v.state := S_WP_SPECIAL_REQUEST_BUSIF_ONLY;
                        end if;
                        if (wpai.gnt_busif = '1' and wpbifi.busif_busy = '0') then
                            v.state := S_WP_SPECIAL;
                        end if;
                    elsif (wpi.port_rlink_wcond = '1') then
                        -- Link current address (LL operation)...
                        v.link_adr := wpi.port_adr;
                        v.link_valid := '1';
                    end if;
                -- Additional state for direct memory access...
                when S_WP_DIRECT =>
                    -- Issue "direct write" operation...
                    vwpao.req_busif := '1';
                    vwpbifo.busif_op := BIO_DIRECT_WRITE;
                    if (wpbifi.busif_busy = '1') then
                        -- Now the BUSIF is busy and has captured the data => can ack and complete
                        vwpo.port_ack := '1';
                        v.state := S_WP_INIT;
                    end if;
                -- Additional states for normal access...
                when S_WP_REQUEST_LINELOCK_ONLY =>
                    -- We got a grant for 'tagr', but not the 'linelock'
                    -- => We must release everything except the 'linelock' to avoid a deadlock
                    vwpao.req_linelock := '1';
                    if (wpai.gnt_linelock = '1') then v.state := S_WP_INIT; end if;
                when S_WP_READ_TAG =>
                    -- Capture the tag and request the bank...
                    vwpao.req_linelock := '1';
                    if (wpi.port_bsel /= X"F") then bank_req_rd := '1'; end if;
                    vwpco.tag_out := wpci.tag_in; -- for bank reading to output the correct cache way
                    v.tag := wpci.tag_in;
                    if (wpci.tag_in.valid = '1') then
                        if (CFG_NUT_HISTOGRAM) then
                            if (r.hist_miss = '0') then
                                hist_cache_write_miss.abort <= '1';
                            end if;
                        end if;
                        -- Cache hit...
                        if (wpi.port_bsel = X"F") then
                            if (wpci.tag_in.dirty = '1') then
                                v.state := S_WP_WRITE_BANK;
                            else
                                v.state := S_WP_WRITE_TAG1_AND_BANK;
                            end if;
                        elsif (bank_gnt = '1') then
                            v.state := S_WP_READ_BANK;
                        else
                            v.state := S_WP_HAVE_TAG_REQUEST_BANK;
                        end if;
                    else
                        if (CFG_NUT_HISTOGRAM) then
                            v.hist_miss := '1';
                        end if;
                        hist_cache_write_hit.abort <= '1';
                        v.state := S_WP_MISS;
                    end if;
                when S_WP_HAVE_TAG_REQUEST_BANK =>
                    vwpao.req_linelock := '1';
                    bank_req_rd := '1';
                    if (bank_gnt = '1') then v.state := S_WP_READ_BANK; end if;
                when S_WP_READ_BANK =>
                    -- read old word (for part-word write only)...
                    vwpao.req_linelock := '1';
                    bank_req_rd := '1';
                    v.data := wpci.bank_data_in;
                    if (r.tag.dirty = '1') then v.state := S_WP_WRITE_BANK;
                    else v.state := S_WP_WRITE_TAG1_AND_BANK;
                    end if;
                when S_WP_WRITE_TAG1_AND_BANK =>
                    vwpao.req_linelock := '1';
                    vwpao.req_tagw := '1';
                    vwpco.tag_out.dirty := '1';
                    bank_req_rd := '1';
                    --vwpco.bank_data_out := combine_data(wpi.port_bsel, r.data, wpi.port_data);
                    if (bank_gnt = '1') then
                        vwpco.bank_wr := '1';
                        v.state := S_WP_WRITE_TAG1;
                    end if;
                    if (wpai.gnt_tagw = '1') then
                        vwpco.tag_wr := '1';
                        v.state := S_WP_WRITE_TAG2_AND_BANK;
                    end if;
                    if (bank_gnt = '1' and wpai.gnt_tagw = '1') then
                        v.state := S_WP_WRITE_TAG2;
                    end if;
                when S_WP_WRITE_TAG2_AND_BANK =>
                    vwpao.req_linelock := '1';
                    vwpao.req_tagw := '1';
                    vwpco.tag_wr := '1';
                    vwpco.tag_out.dirty := '1';
                    bank_req_rd := '1';
                    --vwpco.bank_data_out := combine_data(wpi.port_bsel, r.data, wpi.port_data);
                    if (bank_gnt = '1') then
                        hist_cache_write_hit.stop <= '1';
                        hist_cache_write_miss.stop <= '1';
                        vwpao.req_linelock := '0';
                        vwpco.bank_wr := '1';
                        vwpo.port_ack := '1'; -- can acknowledge to port now (write to bank and tag must be commited!)
                        v.state := S_WP_INIT;
                    else
                        v.state := S_WP_WRITE_BANK;
                    end if;
                when S_WP_WRITE_TAG1 =>
                    vwpao.req_linelock := '1';
                    vwpao.req_tagw := '1';
                    vwpco.tag_out.dirty := '1';
                    if (wpai.gnt_tagw = '1') then
                        vwpco.tag_wr := '1';
                        v.state := S_WP_WRITE_TAG2;
                    end if;
                when S_WP_WRITE_TAG2 =>
                    hist_cache_write_hit.stop <= '1';
                    hist_cache_write_miss.stop <= '1';
                    vwpao.req_linelock := '0';
                    vwpao.req_tagw := '1';
                    vwpco.tag_out.dirty := '1';
                    vwpco.tag_wr := '1';
                    vwpo.port_ack := '1'; -- can acknowledge to port now (write to bank and tag must be commited!)
                    v.state := S_WP_INIT;
                when S_WP_WRITE_BANK =>
                    vwpao.req_linelock := '1';
                    bank_req_rd := '1';
                    --vwpco.bank_data_out := combine_data(wpi.port_bsel, r.data, wpi.port_data);
                    if (bank_gnt = '1') then
                        hist_cache_write_hit.stop <= '1';
                        hist_cache_write_miss.stop <= '1';
                        vwpao.req_linelock := '0';
                        vwpco.bank_wr := '1';
                        vwpo.port_ack := '1'; -- can acknowledge to port now (write to bank must be commited!)
                        v.state := S_WP_INIT;
                    end if;
                    -- Can we accept a new request already in this state?
                    -- -> No, 'tagr' must not be requested while bank is held (deadlock)

                    -- The following states handle a cache miss & replace a cache line.
                when S_WP_MISS =>
                -- Entry state for a cache miss. First, we must request and acquire the BusIf and potentially re-acquire the line lock...
                    vwpao.req_busif := '1';
                    vwpao.req_linelock := '1';
                    if (wpai.gnt_busif = '1' and wpbifi.busif_busy = '0' and wpai.gnt_linelock = '1') then
                        v.state := S_WP_RECHECK;
                    elsif (wpai.gnt_busif = '0' and wpai.gnt_linelock = '1') then
                        v.state := S_WP_REQUEST_BUSIF_ONLY;
                    end if;
                when S_WP_REQUEST_BUSIF_ONLY =>
                    -- Release the line lock and request the BusIf only to avoid deadlocks.
                    vwpao.req_busif := '1';
                    if (wpai.gnt_busif = '1') then v.state := S_WP_MISS; end if;
                when S_WP_RECHECK =>
                    -- Now we have the BusIf and the line lock, and the BusIf
                    -- is idle. We must re-check if there is a cache hit now,
                    -- since some other port may have replaced the cache line in
                    -- between.
                    vwpao.req_busif := '1';
                    vwpao.req_linelock := '1';
                    vwpao.req_tagr := '1';
                    if (wpai.gnt_tagr = '1') then
                        vwpco.tag_rd := '1';
                        v.state := S_WP_RECHECK_READ_TAG;
                    end if;
                when S_WP_RECHECK_READ_TAG =>
                    -- Capture the tag and check it for a cache hit.
                    vwpao.req_busif := '1';
                    vwpao.req_linelock := '1';
                    v.tag := wpci.tag_in;
                    if (wpci.tag_in.valid = '1') then
                        if (wpi.port_bsel = X"F") then
                            if (wpci.tag_in.dirty = '1') then v.state := S_WP_WRITE_BANK;
                            else v.state := S_WP_WRITE_TAG1_AND_BANK;
                            end if;
                        else
                            v.state := S_WP_HAVE_TAG_REQUEST_BANK;
                        end if;
                    else
                        v.state := S_WP_REPLACE;
                    end if;
                when S_WP_REPLACE =>
                    -- Start the replacement by the BusIf.
                    vwpao.req_busif := '1';
                    vwpao.req_linelock := '1';
                    vwpbifo.busif_op := BIO_REPLACE;
                    if (wpbifi.busif_busy = '1') then v.state := S_WP_REPLACE_WAIT_BUSIF; end if;
                when S_WP_REPLACE_WAIT_BUSIF =>
                    -- Wait for the BusIf to complete the replacement.
                    vwpao.req_busif := '1';
                    vwpao.req_linelock := '1';
                    if (wpbifi.busif_busy = '0') then
                        vwpao.req_tagr := '1';
                        if (wpai.gnt_tagr = '1') then
                            vwpco.tag_rd := '1';
                            v.state := S_WP_READ_TAG;
                        else
                            v.state := S_WP_INIT;
                        end if;
                    end if;
                -- States for special operations...
                when S_WP_SPECIAL_REQUEST_BUSIF_ONLY =>
                    vwpao.req_busif := '1';
                    if (wpai.gnt_busif = '1') then v.state := S_WP_INIT; end if;
                when S_WP_SPECIAL =>
                    vwpao.req_busif := '1';
                    vwpao.req_linelock := '1';
                    if (wpi.port_writeback = '1' and wpi.port_invalidate = '1') then 
                        vwpbifo.busif_op := BIO_FLUSH;
                    elsif (wpi.port_writeback = '1') then
                        vwpbifo.busif_op := BIO_WRITEBACK;
                    else
                        vwpbifo.busif_op := BIO_INVALIDATE;
                    end if;
                    if (wpbifi.busif_busy = '1') then
                        v.state := S_WP_SPECIAL_WAIT_COMPLETE;
                    end if;
                when S_WP_SPECIAL_WAIT_COMPLETE =>
                    vwpao.req_busif := '1';
                    vwpao.req_linelock := '1';
                    if (wpbifi.busif_busy = '0') then
                        -- The BusIf has completed -> can ack and complete
                        vwpao.req_linelock := '0';
                        vwpo.port_ack := '1';
                        v.state := S_WP_INIT;
                    end if;
                when others =>
                    v.state := S_WP_INIT;
            end case;
        end if;

        -- Set derived outputs...
        vwpao.req_bank(conv_integer(bank)) := bank_req_rd;
        vwpco.bank_rd := bank_req_rd;

        wpao <= vwpao;
        wpco <= vwpco;
        wpo <= vwpo;
        wpbifo <= vwpbifo;

        rin <= v;

    end process;

    regs : process (clk)
    begin
        if (clk'event and clk = '1') then
            r <= rin;
        end if;
    end process;

end rtl;
