--------------------------------------------------------------------------------
-- This file is part of the ParaNut project.
-- 
-- Copyright (C) 2013  Michael Seider, Hochschule Augsburg
-- michael.seider@hs-augsburg.de
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
-- Description:
--  Readport module for the MEMU.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library paranut;
use paranut.paranut_config.all;
use paranut.types.all;
use paranut.memu_lib.all;
use paranut.paranut_lib.all;
use paranut.histogram.all;

entity mreadport is
        port (
                 clk    : in std_logic;
                 reset  : in std_logic;
                 -- With (CPU) port...
                 rpi    : in readport_in_type;
                 rpo    : out readport_out_type;
                 -- With cache...
                 rpci   : in readport_cache_in_type;
                 rpco   : out readport_cache_out_type;
                 -- With BUSIF...
                 rpbifi : in readport_busif_in_type;
                 rpbifo : out readport_busif_out_type;
                 -- Request & grant lines...
                 rpai   : in readport_arbiter_in_type;
                 rpao   : out readport_arbiter_out_type;
                 -- Histogram...
                 hist_cache_read_hit  : out hist_ctrl_type;
                 hist_cache_read_miss : out hist_ctrl_type
             );
end mreadport;

architecture rtl of mreadport is
    -- - Address information for tag is routed around this module from 'port_adr', for bank from 'port_adr' AND 'way_out'.

    -- - All input ports must be held until 'port_ack' is asserted, at least for one cycle.
    -- - 'port_ack' is issued for exactly one cycle (no full handshake).
    -- - 'port_ack' is issued one cycle before the data is valid (pipelining).
    -- - The next request may be issued at earliest one cycle after 'port_ack' was asserted (which is the same cycle the data is delivered).
    -- - ('port_ack' may be asserted already in the same cycle as the request was issued.) -> minumum latency on cache hit is presently 2 clocks
    -- - If 'port_direct' is set, nothing happens with the cache (i.e. no invalidation).
    --   Hence, 'port_direct' = 0/1 should not be mixed for one address.
    -- - On a 'busif_hit' the next state must set "vrpo.port_data = rpbifi.busif_data" (which is the default for all states)

    type state_type is (S_RP_INIT, S_RP_DIRECT_WAIT_BUSIF,
    S_RP_REQUEST_TAG_ONLY, S_RP_READ_TAG, S_RP_READ_BANK, S_RP_MISS_WAIT_BUSIF,
    S_RP_MISS_REQUEST_TAG, S_RP_MISS_READ_TAG, S_RP_MISS_REPLACE);

    type registers is record
        state    : state_type;
        bank_sel : std_logic_vector(CFG_MEMU_CACHE_BANKS_LD-1 downto 0);
    end record;

    signal r, rin : registers;

begin

    comb : process (r, reset, rpi, rpci, rpbifi, rpai)
        variable v : registers;
        -- Output variables
        variable vrpo    : readport_out_type;
        variable vrpbifo : readport_busif_out_type;
        variable vrpco   : readport_cache_out_type;
        variable vrpao   : readport_arbiter_out_type;
        -- Helper variables...
        variable busif_hit          : std_logic;
        variable index              : std_logic_vector(CFG_MEMU_CACHE_SETS_LD-1 downto 0);
        variable bank               : std_logic_vector(CFG_MEMU_CACHE_BANKS_LD-1 downto 0);
        variable bank_req_rd        : std_logic;
        variable tagr_gnt, bank_gnt : std_logic;
    begin

        v := r;

        hist_cache_read_hit.start <= '0';
        hist_cache_read_hit.stop <= '0';
        hist_cache_read_hit.abort <= '0';
        hist_cache_read_miss.start <= '0';
        hist_cache_read_miss.stop <= '0';
        hist_cache_read_miss.abort <= '0';

        -- Default for outputs...
        vrpo.port_ack := '0';
        vrpo.port_data := rpbifi.busif_data;

        vrpao.req_busif := '0';
        vrpao.req_tagr := '0';
        vrpao.req_bank := (others => '0');

        vrpbifo.busif_op := BIO_NOTHING;

        vrpco.tag_rd := '0';
        vrpco.bank_sel := r.bank_sel;
        vrpco.way_out := rpci.tag_in.way; --TODO: need a register for this?

        -- Helper variables...
        busif_hit := rpbifi.busif_data_valid(conv_integer(rpi.port_adr(BANK_OF_ADDR_RANGE)))
        and conv_std_logic(rpi.port_adr(31 downto 2) = rpbifi.busif_adr(31 downto 2));
        index := rpi.port_adr(INDEX_OF_ADDR_RANGE);
        bank := rpi.port_adr(BANK_OF_ADDR_RANGE);
        bank_req_rd := '0';
        tagr_gnt := rpai.gnt_tagr;
        bank_gnt := rpai.gnt_bank(conv_integer(bank));
        
        if (reset = '1') then
            v.state := S_RP_INIT;
        else
            case r.state is
                when S_RP_INIT =>
                    -- Initial state: On new request, initiate all actions for the first cycle
                    if (rpi.port_rd = '1') then
                        if (rpi.port_direct = '1') then
                            -- uncached memory access...
                            vrpbifo.busif_op := BIO_DIRECT_READ;
                            vrpao.req_busif := '1';
                            if (rpai.gnt_busif = '1') then v.state := S_RP_DIRECT_WAIT_BUSIF; end if;
                        else
                            hist_cache_read_hit.start <= '1';
                            hist_cache_read_miss.start <= '1';
                            -- cached memory access...
                            if (busif_hit = '1') then
                                hist_cache_read_hit.abort <= '1';
                                hist_cache_read_miss.abort <= '1';
                                vrpo.port_ack := '1';
                            else
                                vrpao.req_tagr := '1';
                                if (tagr_gnt = '1') then
                                    vrpco.tag_rd := '1';
                                    v.state := S_RP_READ_TAG;
                                end if;
                            end if;
                        end if;
                    end if;
                when S_RP_DIRECT_WAIT_BUSIF =>
                    -- Direct access: Wait for response from BUSIF
                    vrpbifo.busif_op := BIO_DIRECT_READ;
                    vrpao.req_busif := '1';
                    if (busif_hit = '1') then
                        vrpo.port_ack := '1';
                        v.state := S_RP_INIT;
                    end if;
                when S_RP_READ_TAG =>
                    -- Capture the tag (which was granted last state)
                    -- keep req_tagr to hold tag output
                    vrpao.req_tagr := '1';
                    if (rpci.tag_in.valid = '1') then
                        hist_cache_read_miss.abort <= '1';
                        -- Cache hit...
                        bank_req_rd := '1';
                        if (bank_gnt = '1') then
                            hist_cache_read_hit.stop <= '1';
                            vrpao.req_tagr := '0';
                            v.bank_sel := bank;
                            vrpo.port_ack := '1';
                            v.state := S_RP_READ_BANK;
                        end if;
                    else
                        hist_cache_read_hit.abort <= '1';
                        v.state := S_RP_MISS_WAIT_BUSIF;
                    end if;
                when S_RP_READ_BANK =>
                    -- Read the bank & complete...
                    vrpo.port_data := rpci.bank_data_in;
                    v.state := S_RP_INIT;

                    -- On new request, initiate all actions for the first cycle
                    if (rpi.port_rd = '1') then
                        if (rpi.port_direct = '1') then
                            -- uncached memory access...
                            vrpbifo.busif_op := BIO_DIRECT_READ;
                            vrpao.req_busif := '1';
                            if (rpai.gnt_busif = '1') then v.state := S_RP_DIRECT_WAIT_BUSIF; end if;
                        else
                            hist_cache_read_hit.start <= '1';
                            hist_cache_read_miss.start <= '1';
                            -- cached memory access...
                            if (busif_hit = '1') then
                                hist_cache_read_hit.abort <= '1';
                                hist_cache_read_miss.abort <= '1';
                                vrpo.port_ack := '1';
                            else
                                vrpao.req_tagr := '1';
                                if (tagr_gnt = '1') then
                                    vrpco.tag_rd := '1';
                                    v.state := S_RP_READ_TAG;
                                end if;
                            end if;
                        end if;
                    end if;
                when S_RP_MISS_WAIT_BUSIF =>
                    -- Cache miss detected: Wait until we get the BusIF and the
                    -- BusIF becomes idle and catch an incidental BusIF hit if it
                    -- happens.
                    vrpao.req_busif := '1';
                    if (busif_hit = '1') then
                        hist_cache_read_miss.stop <= '1';
                        vrpo.port_ack := '1';
                        v.state := S_RP_INIT;
                    elsif (rpai.gnt_busif = '1' and rpbifi.busif_busy = '0') then
                        v.state := S_RP_MISS_REQUEST_TAG;
                    end if;
                when S_RP_MISS_REQUEST_TAG =>
                    -- Request the tag again to check for a cache hit. The BusIF
                    -- might already have replaced the cache line during
                    -- 'S_RP_MISS_WAIT_BUSIF' on the request of some other port,
                    -- and that data may have even been modified by a write port!
                    -- Hence, replacing that cache line again would lead to wrong
                    -- data.
                    vrpao.req_busif := '1';
                    vrpao.req_tagr := '1';
                    if (tagr_gnt = '1') then
                        vrpco.tag_rd := '1';
                        v.state := S_RP_MISS_READ_TAG;
                    end if;
                when S_RP_MISS_READ_TAG =>
                    -- read the tag & check for a cache hit
                    vrpao.req_busif := '1';
                    -- keep req_tagr to hold tag output
                    vrpao.req_tagr := '1';
                    if (rpci.tag_in.valid = '1') then
                        bank_req_rd := '1';
                        if (bank_gnt = '1') then
                            hist_cache_read_miss.stop <= '1';
                            vrpao.req_tagr := '0';
                            v.bank_sel := bank;
                            vrpo.port_ack := '1';
                            v.state := S_RP_READ_BANK;
                        end if;
                    else
                        v.state := S_RP_MISS_REPLACE;
                    end if;
                when S_RP_MISS_REPLACE =>
                    -- Run the replacement and wait for the BusIF hit which MUST come some time
                    vrpao.req_busif := '1';
                    vrpbifo.busif_op := BIO_REPLACE;
                    if (busif_hit = '1') then
                        hist_cache_read_miss.stop <= '1';
                        vrpo.port_ack := '1';
                        v.state := S_RP_INIT;
                    end if;
                when others =>
                    v.state := S_RP_INIT;
            end case;
        end if;

        -- Set derived outputs...
        vrpao.req_bank(conv_integer(bank)) := bank_req_rd;
        vrpco.bank_rd := bank_req_rd;

        rpo <= vrpo;
        rpbifo <= vrpbifo;
        rpco <= vrpco;
        rpao <= vrpao;

        rin <= v;

    end process;

    regs : process (clk)
    begin
        if (clk'event and clk = '1') then
            r <= rin;
        end if;
    end process;

end rtl;
