library ieee;
use ieee.std_logic_1164.all;

library paranut;
use paranut.types.all;

package prog_mem is

	constant PROG_SIZE : integer := 93664;

	constant PROG_DATA : mem_type(0 to PROG_SIZE/4-1) := (
		16#0000# => X"00000000",
		16#0001# => X"00000000",
		16#0002# => X"00000000",
		16#0003# => X"00000000",
		16#0004# => X"00000000",
		16#0005# => X"00000000",
		16#0006# => X"00000000",
		16#0007# => X"00000000",
		16#0008# => X"00000000",
		16#0009# => X"00000000",
		16#000a# => X"00000000",
		16#000b# => X"00000000",
		16#000c# => X"00000000",
		16#000d# => X"00000000",
		16#000e# => X"00000000",
		16#000f# => X"00000000",
		16#0010# => X"00000000",
		16#0011# => X"00000000",
		16#0012# => X"00000000",
		16#0013# => X"00000000",
		16#0014# => X"00000000",
		16#0015# => X"00000000",
		16#0016# => X"00000000",
		16#0017# => X"00000000",
		16#0018# => X"00000000",
		16#0019# => X"00000000",
		16#001a# => X"00000000",
		16#001b# => X"00000000",
		16#001c# => X"00000000",
		16#001d# => X"00000000",
		16#001e# => X"00000000",
		16#001f# => X"00000000",
		16#0020# => X"00000000",
		16#0021# => X"00000000",
		16#0022# => X"00000000",
		16#0023# => X"00000000",
		16#0024# => X"00000000",
		16#0025# => X"00000000",
		16#0026# => X"00000000",
		16#0027# => X"00000000",
		16#0028# => X"00000000",
		16#0029# => X"00000000",
		16#002a# => X"00000000",
		16#002b# => X"00000000",
		16#002c# => X"00000000",
		16#002d# => X"00000000",
		16#002e# => X"00000000",
		16#002f# => X"00000000",
		16#0030# => X"00000000",
		16#0031# => X"00000000",
		16#0032# => X"00000000",
		16#0033# => X"00000000",
		16#0034# => X"00000000",
		16#0035# => X"00000000",
		16#0036# => X"00000000",
		16#0037# => X"00000000",
		16#0038# => X"00000000",
		16#0039# => X"00000000",
		16#003a# => X"00000000",
		16#003b# => X"00000000",
		16#003c# => X"00000000",
		16#003d# => X"00000000",
		16#003e# => X"00000000",
		16#003f# => X"00000000",
		16#0040# => X"18000000",
		16#0041# => X"18200000",
		16#0042# => X"18400000",
		16#0043# => X"18600000",
		16#0044# => X"18800000",
		16#0045# => X"18a00000",
		16#0046# => X"18c00000",
		16#0047# => X"18e00000",
		16#0048# => X"19000000",
		16#0049# => X"19200000",
		16#004a# => X"19400000",
		16#004b# => X"19600000",
		16#004c# => X"19800000",
		16#004d# => X"19a00000",
		16#004e# => X"19c00000",
		16#004f# => X"19e00000",
		16#0050# => X"1a000000",
		16#0051# => X"1a200000",
		16#0052# => X"1a400000",
		16#0053# => X"1a600000",
		16#0054# => X"1a800000",
		16#0055# => X"1aa00000",
		16#0056# => X"1ac00000",
		16#0057# => X"1ae00000",
		16#0058# => X"1b000000",
		16#0059# => X"1b200000",
		16#005a# => X"1b400000",
		16#005b# => X"1b600000",
		16#005c# => X"1b800000",
		16#005d# => X"1ba00000",
		16#005e# => X"1bc00000",
		16#005f# => X"1be00000",
		16#0060# => X"a8200001",
		16#0061# => X"c0000811",
		16#0062# => X"c1400000",
		16#0063# => X"18800000",
		16#0064# => X"a8842028",
		16#0065# => X"44002000",
		16#0066# => X"15000000",
		16#0067# => X"00000000",
		16#0068# => X"00000000",
		16#0069# => X"00000000",
		16#006a# => X"00000000",
		16#006b# => X"00000000",
		16#006c# => X"00000000",
		16#006d# => X"00000000",
		16#006e# => X"00000000",
		16#006f# => X"00000000",
		16#0070# => X"00000000",
		16#0071# => X"00000000",
		16#0072# => X"00000000",
		16#0073# => X"00000000",
		16#0074# => X"00000000",
		16#0075# => X"00000000",
		16#0076# => X"00000000",
		16#0077# => X"00000000",
		16#0078# => X"00000000",
		16#0079# => X"00000000",
		16#007a# => X"00000000",
		16#007b# => X"00000000",
		16#007c# => X"00000000",
		16#007d# => X"00000000",
		16#007e# => X"00000000",
		16#007f# => X"00000000",
		16#0080# => X"9c21ff00",
		16#0081# => X"d4011804",
		16#0082# => X"d4012008",
		16#0083# => X"b4600010",
		16#0084# => X"000020f4",
		16#0085# => X"b4800020",
		16#0086# => X"00000000",
		16#0087# => X"00000000",
		16#0088# => X"00000000",
		16#0089# => X"00000000",
		16#008a# => X"00000000",
		16#008b# => X"00000000",
		16#008c# => X"00000000",
		16#008d# => X"00000000",
		16#008e# => X"00000000",
		16#008f# => X"00000000",
		16#0090# => X"00000000",
		16#0091# => X"00000000",
		16#0092# => X"00000000",
		16#0093# => X"00000000",
		16#0094# => X"00000000",
		16#0095# => X"00000000",
		16#0096# => X"00000000",
		16#0097# => X"00000000",
		16#0098# => X"00000000",
		16#0099# => X"00000000",
		16#009a# => X"00000000",
		16#009b# => X"00000000",
		16#009c# => X"00000000",
		16#009d# => X"00000000",
		16#009e# => X"00000000",
		16#009f# => X"00000000",
		16#00a0# => X"00000000",
		16#00a1# => X"00000000",
		16#00a2# => X"00000000",
		16#00a3# => X"00000000",
		16#00a4# => X"00000000",
		16#00a5# => X"00000000",
		16#00a6# => X"00000000",
		16#00a7# => X"00000000",
		16#00a8# => X"00000000",
		16#00a9# => X"00000000",
		16#00aa# => X"00000000",
		16#00ab# => X"00000000",
		16#00ac# => X"00000000",
		16#00ad# => X"00000000",
		16#00ae# => X"00000000",
		16#00af# => X"00000000",
		16#00b0# => X"00000000",
		16#00b1# => X"00000000",
		16#00b2# => X"00000000",
		16#00b3# => X"00000000",
		16#00b4# => X"00000000",
		16#00b5# => X"00000000",
		16#00b6# => X"00000000",
		16#00b7# => X"00000000",
		16#00b8# => X"00000000",
		16#00b9# => X"00000000",
		16#00ba# => X"00000000",
		16#00bb# => X"00000000",
		16#00bc# => X"00000000",
		16#00bd# => X"00000000",
		16#00be# => X"00000000",
		16#00bf# => X"00000000",
		16#00c0# => X"9c21ff00",
		16#00c1# => X"d4011804",
		16#00c2# => X"d4012008",
		16#00c3# => X"b4600010",
		16#00c4# => X"000020b4",
		16#00c5# => X"b4800020",
		16#00c6# => X"00000000",
		16#00c7# => X"00000000",
		16#00c8# => X"00000000",
		16#00c9# => X"00000000",
		16#00ca# => X"00000000",
		16#00cb# => X"00000000",
		16#00cc# => X"00000000",
		16#00cd# => X"00000000",
		16#00ce# => X"00000000",
		16#00cf# => X"00000000",
		16#00d0# => X"00000000",
		16#00d1# => X"00000000",
		16#00d2# => X"00000000",
		16#00d3# => X"00000000",
		16#00d4# => X"00000000",
		16#00d5# => X"00000000",
		16#00d6# => X"00000000",
		16#00d7# => X"00000000",
		16#00d8# => X"00000000",
		16#00d9# => X"00000000",
		16#00da# => X"00000000",
		16#00db# => X"00000000",
		16#00dc# => X"00000000",
		16#00dd# => X"00000000",
		16#00de# => X"00000000",
		16#00df# => X"00000000",
		16#00e0# => X"00000000",
		16#00e1# => X"00000000",
		16#00e2# => X"00000000",
		16#00e3# => X"00000000",
		16#00e4# => X"00000000",
		16#00e5# => X"00000000",
		16#00e6# => X"00000000",
		16#00e7# => X"00000000",
		16#00e8# => X"00000000",
		16#00e9# => X"00000000",
		16#00ea# => X"00000000",
		16#00eb# => X"00000000",
		16#00ec# => X"00000000",
		16#00ed# => X"00000000",
		16#00ee# => X"00000000",
		16#00ef# => X"00000000",
		16#00f0# => X"00000000",
		16#00f1# => X"00000000",
		16#00f2# => X"00000000",
		16#00f3# => X"00000000",
		16#00f4# => X"00000000",
		16#00f5# => X"00000000",
		16#00f6# => X"00000000",
		16#00f7# => X"00000000",
		16#00f8# => X"00000000",
		16#00f9# => X"00000000",
		16#00fa# => X"00000000",
		16#00fb# => X"00000000",
		16#00fc# => X"00000000",
		16#00fd# => X"00000000",
		16#00fe# => X"00000000",
		16#00ff# => X"00000000",
		16#0100# => X"9c21ff00",
		16#0101# => X"d4011804",
		16#0102# => X"d4012008",
		16#0103# => X"b4600010",
		16#0104# => X"00002074",
		16#0105# => X"b4800020",
		16#0106# => X"00000000",
		16#0107# => X"00000000",
		16#0108# => X"00000000",
		16#0109# => X"00000000",
		16#010a# => X"00000000",
		16#010b# => X"00000000",
		16#010c# => X"00000000",
		16#010d# => X"00000000",
		16#010e# => X"00000000",
		16#010f# => X"00000000",
		16#0110# => X"00000000",
		16#0111# => X"00000000",
		16#0112# => X"00000000",
		16#0113# => X"00000000",
		16#0114# => X"00000000",
		16#0115# => X"00000000",
		16#0116# => X"00000000",
		16#0117# => X"00000000",
		16#0118# => X"00000000",
		16#0119# => X"00000000",
		16#011a# => X"00000000",
		16#011b# => X"00000000",
		16#011c# => X"00000000",
		16#011d# => X"00000000",
		16#011e# => X"00000000",
		16#011f# => X"00000000",
		16#0120# => X"00000000",
		16#0121# => X"00000000",
		16#0122# => X"00000000",
		16#0123# => X"00000000",
		16#0124# => X"00000000",
		16#0125# => X"00000000",
		16#0126# => X"00000000",
		16#0127# => X"00000000",
		16#0128# => X"00000000",
		16#0129# => X"00000000",
		16#012a# => X"00000000",
		16#012b# => X"00000000",
		16#012c# => X"00000000",
		16#012d# => X"00000000",
		16#012e# => X"00000000",
		16#012f# => X"00000000",
		16#0130# => X"00000000",
		16#0131# => X"00000000",
		16#0132# => X"00000000",
		16#0133# => X"00000000",
		16#0134# => X"00000000",
		16#0135# => X"00000000",
		16#0136# => X"00000000",
		16#0137# => X"00000000",
		16#0138# => X"00000000",
		16#0139# => X"00000000",
		16#013a# => X"00000000",
		16#013b# => X"00000000",
		16#013c# => X"00000000",
		16#013d# => X"00000000",
		16#013e# => X"00000000",
		16#013f# => X"00000000",
		16#0140# => X"9c21ff00",
		16#0141# => X"d4011804",
		16#0142# => X"d4012008",
		16#0143# => X"b4600010",
		16#0144# => X"00002034",
		16#0145# => X"b4800020",
		16#0146# => X"00000000",
		16#0147# => X"00000000",
		16#0148# => X"00000000",
		16#0149# => X"00000000",
		16#014a# => X"00000000",
		16#014b# => X"00000000",
		16#014c# => X"00000000",
		16#014d# => X"00000000",
		16#014e# => X"00000000",
		16#014f# => X"00000000",
		16#0150# => X"00000000",
		16#0151# => X"00000000",
		16#0152# => X"00000000",
		16#0153# => X"00000000",
		16#0154# => X"00000000",
		16#0155# => X"00000000",
		16#0156# => X"00000000",
		16#0157# => X"00000000",
		16#0158# => X"00000000",
		16#0159# => X"00000000",
		16#015a# => X"00000000",
		16#015b# => X"00000000",
		16#015c# => X"00000000",
		16#015d# => X"00000000",
		16#015e# => X"00000000",
		16#015f# => X"00000000",
		16#0160# => X"00000000",
		16#0161# => X"00000000",
		16#0162# => X"00000000",
		16#0163# => X"00000000",
		16#0164# => X"00000000",
		16#0165# => X"00000000",
		16#0166# => X"00000000",
		16#0167# => X"00000000",
		16#0168# => X"00000000",
		16#0169# => X"00000000",
		16#016a# => X"00000000",
		16#016b# => X"00000000",
		16#016c# => X"00000000",
		16#016d# => X"00000000",
		16#016e# => X"00000000",
		16#016f# => X"00000000",
		16#0170# => X"00000000",
		16#0171# => X"00000000",
		16#0172# => X"00000000",
		16#0173# => X"00000000",
		16#0174# => X"00000000",
		16#0175# => X"00000000",
		16#0176# => X"00000000",
		16#0177# => X"00000000",
		16#0178# => X"00000000",
		16#0179# => X"00000000",
		16#017a# => X"00000000",
		16#017b# => X"00000000",
		16#017c# => X"00000000",
		16#017d# => X"00000000",
		16#017e# => X"00000000",
		16#017f# => X"00000000",
		16#0180# => X"9c21ff00",
		16#0181# => X"d4011804",
		16#0182# => X"d4012008",
		16#0183# => X"b4600010",
		16#0184# => X"00001ff4",
		16#0185# => X"b4800020",
		16#0186# => X"00000000",
		16#0187# => X"00000000",
		16#0188# => X"00000000",
		16#0189# => X"00000000",
		16#018a# => X"00000000",
		16#018b# => X"00000000",
		16#018c# => X"00000000",
		16#018d# => X"00000000",
		16#018e# => X"00000000",
		16#018f# => X"00000000",
		16#0190# => X"00000000",
		16#0191# => X"00000000",
		16#0192# => X"00000000",
		16#0193# => X"00000000",
		16#0194# => X"00000000",
		16#0195# => X"00000000",
		16#0196# => X"00000000",
		16#0197# => X"00000000",
		16#0198# => X"00000000",
		16#0199# => X"00000000",
		16#019a# => X"00000000",
		16#019b# => X"00000000",
		16#019c# => X"00000000",
		16#019d# => X"00000000",
		16#019e# => X"00000000",
		16#019f# => X"00000000",
		16#01a0# => X"00000000",
		16#01a1# => X"00000000",
		16#01a2# => X"00000000",
		16#01a3# => X"00000000",
		16#01a4# => X"00000000",
		16#01a5# => X"00000000",
		16#01a6# => X"00000000",
		16#01a7# => X"00000000",
		16#01a8# => X"00000000",
		16#01a9# => X"00000000",
		16#01aa# => X"00000000",
		16#01ab# => X"00000000",
		16#01ac# => X"00000000",
		16#01ad# => X"00000000",
		16#01ae# => X"00000000",
		16#01af# => X"00000000",
		16#01b0# => X"00000000",
		16#01b1# => X"00000000",
		16#01b2# => X"00000000",
		16#01b3# => X"00000000",
		16#01b4# => X"00000000",
		16#01b5# => X"00000000",
		16#01b6# => X"00000000",
		16#01b7# => X"00000000",
		16#01b8# => X"00000000",
		16#01b9# => X"00000000",
		16#01ba# => X"00000000",
		16#01bb# => X"00000000",
		16#01bc# => X"00000000",
		16#01bd# => X"00000000",
		16#01be# => X"00000000",
		16#01bf# => X"00000000",
		16#01c0# => X"9c21ff00",
		16#01c1# => X"d4011804",
		16#01c2# => X"d4012008",
		16#01c3# => X"b4600010",
		16#01c4# => X"00001fb4",
		16#01c5# => X"b4800020",
		16#01c6# => X"00000000",
		16#01c7# => X"00000000",
		16#01c8# => X"00000000",
		16#01c9# => X"00000000",
		16#01ca# => X"00000000",
		16#01cb# => X"00000000",
		16#01cc# => X"00000000",
		16#01cd# => X"00000000",
		16#01ce# => X"00000000",
		16#01cf# => X"00000000",
		16#01d0# => X"00000000",
		16#01d1# => X"00000000",
		16#01d2# => X"00000000",
		16#01d3# => X"00000000",
		16#01d4# => X"00000000",
		16#01d5# => X"00000000",
		16#01d6# => X"00000000",
		16#01d7# => X"00000000",
		16#01d8# => X"00000000",
		16#01d9# => X"00000000",
		16#01da# => X"00000000",
		16#01db# => X"00000000",
		16#01dc# => X"00000000",
		16#01dd# => X"00000000",
		16#01de# => X"00000000",
		16#01df# => X"00000000",
		16#01e0# => X"00000000",
		16#01e1# => X"00000000",
		16#01e2# => X"00000000",
		16#01e3# => X"00000000",
		16#01e4# => X"00000000",
		16#01e5# => X"00000000",
		16#01e6# => X"00000000",
		16#01e7# => X"00000000",
		16#01e8# => X"00000000",
		16#01e9# => X"00000000",
		16#01ea# => X"00000000",
		16#01eb# => X"00000000",
		16#01ec# => X"00000000",
		16#01ed# => X"00000000",
		16#01ee# => X"00000000",
		16#01ef# => X"00000000",
		16#01f0# => X"00000000",
		16#01f1# => X"00000000",
		16#01f2# => X"00000000",
		16#01f3# => X"00000000",
		16#01f4# => X"00000000",
		16#01f5# => X"00000000",
		16#01f6# => X"00000000",
		16#01f7# => X"00000000",
		16#01f8# => X"00000000",
		16#01f9# => X"00000000",
		16#01fa# => X"00000000",
		16#01fb# => X"00000000",
		16#01fc# => X"00000000",
		16#01fd# => X"00000000",
		16#01fe# => X"00000000",
		16#01ff# => X"00000000",
		16#0200# => X"9c21ff00",
		16#0201# => X"d4011804",
		16#0202# => X"d4012008",
		16#0203# => X"b4600010",
		16#0204# => X"00001f74",
		16#0205# => X"b4800020",
		16#0206# => X"00000000",
		16#0207# => X"00000000",
		16#0208# => X"00000000",
		16#0209# => X"00000000",
		16#020a# => X"00000000",
		16#020b# => X"00000000",
		16#020c# => X"00000000",
		16#020d# => X"00000000",
		16#020e# => X"00000000",
		16#020f# => X"00000000",
		16#0210# => X"00000000",
		16#0211# => X"00000000",
		16#0212# => X"00000000",
		16#0213# => X"00000000",
		16#0214# => X"00000000",
		16#0215# => X"00000000",
		16#0216# => X"00000000",
		16#0217# => X"00000000",
		16#0218# => X"00000000",
		16#0219# => X"00000000",
		16#021a# => X"00000000",
		16#021b# => X"00000000",
		16#021c# => X"00000000",
		16#021d# => X"00000000",
		16#021e# => X"00000000",
		16#021f# => X"00000000",
		16#0220# => X"00000000",
		16#0221# => X"00000000",
		16#0222# => X"00000000",
		16#0223# => X"00000000",
		16#0224# => X"00000000",
		16#0225# => X"00000000",
		16#0226# => X"00000000",
		16#0227# => X"00000000",
		16#0228# => X"00000000",
		16#0229# => X"00000000",
		16#022a# => X"00000000",
		16#022b# => X"00000000",
		16#022c# => X"00000000",
		16#022d# => X"00000000",
		16#022e# => X"00000000",
		16#022f# => X"00000000",
		16#0230# => X"00000000",
		16#0231# => X"00000000",
		16#0232# => X"00000000",
		16#0233# => X"00000000",
		16#0234# => X"00000000",
		16#0235# => X"00000000",
		16#0236# => X"00000000",
		16#0237# => X"00000000",
		16#0238# => X"00000000",
		16#0239# => X"00000000",
		16#023a# => X"00000000",
		16#023b# => X"00000000",
		16#023c# => X"00000000",
		16#023d# => X"00000000",
		16#023e# => X"00000000",
		16#023f# => X"00000000",
		16#0240# => X"9c21ff00",
		16#0241# => X"d4011804",
		16#0242# => X"d4012008",
		16#0243# => X"b4600010",
		16#0244# => X"00001f34",
		16#0245# => X"b4800020",
		16#0246# => X"00000000",
		16#0247# => X"00000000",
		16#0248# => X"00000000",
		16#0249# => X"00000000",
		16#024a# => X"00000000",
		16#024b# => X"00000000",
		16#024c# => X"00000000",
		16#024d# => X"00000000",
		16#024e# => X"00000000",
		16#024f# => X"00000000",
		16#0250# => X"00000000",
		16#0251# => X"00000000",
		16#0252# => X"00000000",
		16#0253# => X"00000000",
		16#0254# => X"00000000",
		16#0255# => X"00000000",
		16#0256# => X"00000000",
		16#0257# => X"00000000",
		16#0258# => X"00000000",
		16#0259# => X"00000000",
		16#025a# => X"00000000",
		16#025b# => X"00000000",
		16#025c# => X"00000000",
		16#025d# => X"00000000",
		16#025e# => X"00000000",
		16#025f# => X"00000000",
		16#0260# => X"00000000",
		16#0261# => X"00000000",
		16#0262# => X"00000000",
		16#0263# => X"00000000",
		16#0264# => X"00000000",
		16#0265# => X"00000000",
		16#0266# => X"00000000",
		16#0267# => X"00000000",
		16#0268# => X"00000000",
		16#0269# => X"00000000",
		16#026a# => X"00000000",
		16#026b# => X"00000000",
		16#026c# => X"00000000",
		16#026d# => X"00000000",
		16#026e# => X"00000000",
		16#026f# => X"00000000",
		16#0270# => X"00000000",
		16#0271# => X"00000000",
		16#0272# => X"00000000",
		16#0273# => X"00000000",
		16#0274# => X"00000000",
		16#0275# => X"00000000",
		16#0276# => X"00000000",
		16#0277# => X"00000000",
		16#0278# => X"00000000",
		16#0279# => X"00000000",
		16#027a# => X"00000000",
		16#027b# => X"00000000",
		16#027c# => X"00000000",
		16#027d# => X"00000000",
		16#027e# => X"00000000",
		16#027f# => X"00000000",
		16#0280# => X"9c21ff00",
		16#0281# => X"d4011804",
		16#0282# => X"d4012008",
		16#0283# => X"b4600010",
		16#0284# => X"00001ef4",
		16#0285# => X"b4800020",
		16#0286# => X"00000000",
		16#0287# => X"00000000",
		16#0288# => X"00000000",
		16#0289# => X"00000000",
		16#028a# => X"00000000",
		16#028b# => X"00000000",
		16#028c# => X"00000000",
		16#028d# => X"00000000",
		16#028e# => X"00000000",
		16#028f# => X"00000000",
		16#0290# => X"00000000",
		16#0291# => X"00000000",
		16#0292# => X"00000000",
		16#0293# => X"00000000",
		16#0294# => X"00000000",
		16#0295# => X"00000000",
		16#0296# => X"00000000",
		16#0297# => X"00000000",
		16#0298# => X"00000000",
		16#0299# => X"00000000",
		16#029a# => X"00000000",
		16#029b# => X"00000000",
		16#029c# => X"00000000",
		16#029d# => X"00000000",
		16#029e# => X"00000000",
		16#029f# => X"00000000",
		16#02a0# => X"00000000",
		16#02a1# => X"00000000",
		16#02a2# => X"00000000",
		16#02a3# => X"00000000",
		16#02a4# => X"00000000",
		16#02a5# => X"00000000",
		16#02a6# => X"00000000",
		16#02a7# => X"00000000",
		16#02a8# => X"00000000",
		16#02a9# => X"00000000",
		16#02aa# => X"00000000",
		16#02ab# => X"00000000",
		16#02ac# => X"00000000",
		16#02ad# => X"00000000",
		16#02ae# => X"00000000",
		16#02af# => X"00000000",
		16#02b0# => X"00000000",
		16#02b1# => X"00000000",
		16#02b2# => X"00000000",
		16#02b3# => X"00000000",
		16#02b4# => X"00000000",
		16#02b5# => X"00000000",
		16#02b6# => X"00000000",
		16#02b7# => X"00000000",
		16#02b8# => X"00000000",
		16#02b9# => X"00000000",
		16#02ba# => X"00000000",
		16#02bb# => X"00000000",
		16#02bc# => X"00000000",
		16#02bd# => X"00000000",
		16#02be# => X"00000000",
		16#02bf# => X"00000000",
		16#02c0# => X"9c21ff00",
		16#02c1# => X"d4011804",
		16#02c2# => X"d4012008",
		16#02c3# => X"b4600010",
		16#02c4# => X"00001eb4",
		16#02c5# => X"b4800020",
		16#02c6# => X"00000000",
		16#02c7# => X"00000000",
		16#02c8# => X"00000000",
		16#02c9# => X"00000000",
		16#02ca# => X"00000000",
		16#02cb# => X"00000000",
		16#02cc# => X"00000000",
		16#02cd# => X"00000000",
		16#02ce# => X"00000000",
		16#02cf# => X"00000000",
		16#02d0# => X"00000000",
		16#02d1# => X"00000000",
		16#02d2# => X"00000000",
		16#02d3# => X"00000000",
		16#02d4# => X"00000000",
		16#02d5# => X"00000000",
		16#02d6# => X"00000000",
		16#02d7# => X"00000000",
		16#02d8# => X"00000000",
		16#02d9# => X"00000000",
		16#02da# => X"00000000",
		16#02db# => X"00000000",
		16#02dc# => X"00000000",
		16#02dd# => X"00000000",
		16#02de# => X"00000000",
		16#02df# => X"00000000",
		16#02e0# => X"00000000",
		16#02e1# => X"00000000",
		16#02e2# => X"00000000",
		16#02e3# => X"00000000",
		16#02e4# => X"00000000",
		16#02e5# => X"00000000",
		16#02e6# => X"00000000",
		16#02e7# => X"00000000",
		16#02e8# => X"00000000",
		16#02e9# => X"00000000",
		16#02ea# => X"00000000",
		16#02eb# => X"00000000",
		16#02ec# => X"00000000",
		16#02ed# => X"00000000",
		16#02ee# => X"00000000",
		16#02ef# => X"00000000",
		16#02f0# => X"00000000",
		16#02f1# => X"00000000",
		16#02f2# => X"00000000",
		16#02f3# => X"00000000",
		16#02f4# => X"00000000",
		16#02f5# => X"00000000",
		16#02f6# => X"00000000",
		16#02f7# => X"00000000",
		16#02f8# => X"00000000",
		16#02f9# => X"00000000",
		16#02fa# => X"00000000",
		16#02fb# => X"00000000",
		16#02fc# => X"00000000",
		16#02fd# => X"00000000",
		16#02fe# => X"00000000",
		16#02ff# => X"00000000",
		16#0300# => X"9c21ff00",
		16#0301# => X"d4011804",
		16#0302# => X"d4012008",
		16#0303# => X"b4600010",
		16#0304# => X"00001e74",
		16#0305# => X"b4800020",
		16#0306# => X"00000000",
		16#0307# => X"00000000",
		16#0308# => X"00000000",
		16#0309# => X"00000000",
		16#030a# => X"00000000",
		16#030b# => X"00000000",
		16#030c# => X"00000000",
		16#030d# => X"00000000",
		16#030e# => X"00000000",
		16#030f# => X"00000000",
		16#0310# => X"00000000",
		16#0311# => X"00000000",
		16#0312# => X"00000000",
		16#0313# => X"00000000",
		16#0314# => X"00000000",
		16#0315# => X"00000000",
		16#0316# => X"00000000",
		16#0317# => X"00000000",
		16#0318# => X"00000000",
		16#0319# => X"00000000",
		16#031a# => X"00000000",
		16#031b# => X"00000000",
		16#031c# => X"00000000",
		16#031d# => X"00000000",
		16#031e# => X"00000000",
		16#031f# => X"00000000",
		16#0320# => X"00000000",
		16#0321# => X"00000000",
		16#0322# => X"00000000",
		16#0323# => X"00000000",
		16#0324# => X"00000000",
		16#0325# => X"00000000",
		16#0326# => X"00000000",
		16#0327# => X"00000000",
		16#0328# => X"00000000",
		16#0329# => X"00000000",
		16#032a# => X"00000000",
		16#032b# => X"00000000",
		16#032c# => X"00000000",
		16#032d# => X"00000000",
		16#032e# => X"00000000",
		16#032f# => X"00000000",
		16#0330# => X"00000000",
		16#0331# => X"00000000",
		16#0332# => X"00000000",
		16#0333# => X"00000000",
		16#0334# => X"00000000",
		16#0335# => X"00000000",
		16#0336# => X"00000000",
		16#0337# => X"00000000",
		16#0338# => X"00000000",
		16#0339# => X"00000000",
		16#033a# => X"00000000",
		16#033b# => X"00000000",
		16#033c# => X"00000000",
		16#033d# => X"00000000",
		16#033e# => X"00000000",
		16#033f# => X"00000000",
		16#0340# => X"9c21ff00",
		16#0341# => X"d4011804",
		16#0342# => X"d4012008",
		16#0343# => X"b4600010",
		16#0344# => X"00001e34",
		16#0345# => X"b4800020",
		16#0346# => X"00000000",
		16#0347# => X"00000000",
		16#0348# => X"00000000",
		16#0349# => X"00000000",
		16#034a# => X"00000000",
		16#034b# => X"00000000",
		16#034c# => X"00000000",
		16#034d# => X"00000000",
		16#034e# => X"00000000",
		16#034f# => X"00000000",
		16#0350# => X"00000000",
		16#0351# => X"00000000",
		16#0352# => X"00000000",
		16#0353# => X"00000000",
		16#0354# => X"00000000",
		16#0355# => X"00000000",
		16#0356# => X"00000000",
		16#0357# => X"00000000",
		16#0358# => X"00000000",
		16#0359# => X"00000000",
		16#035a# => X"00000000",
		16#035b# => X"00000000",
		16#035c# => X"00000000",
		16#035d# => X"00000000",
		16#035e# => X"00000000",
		16#035f# => X"00000000",
		16#0360# => X"00000000",
		16#0361# => X"00000000",
		16#0362# => X"00000000",
		16#0363# => X"00000000",
		16#0364# => X"00000000",
		16#0365# => X"00000000",
		16#0366# => X"00000000",
		16#0367# => X"00000000",
		16#0368# => X"00000000",
		16#0369# => X"00000000",
		16#036a# => X"00000000",
		16#036b# => X"00000000",
		16#036c# => X"00000000",
		16#036d# => X"00000000",
		16#036e# => X"00000000",
		16#036f# => X"00000000",
		16#0370# => X"00000000",
		16#0371# => X"00000000",
		16#0372# => X"00000000",
		16#0373# => X"00000000",
		16#0374# => X"00000000",
		16#0375# => X"00000000",
		16#0376# => X"00000000",
		16#0377# => X"00000000",
		16#0378# => X"00000000",
		16#0379# => X"00000000",
		16#037a# => X"00000000",
		16#037b# => X"00000000",
		16#037c# => X"00000000",
		16#037d# => X"00000000",
		16#037e# => X"00000000",
		16#037f# => X"00000000",
		16#0380# => X"9c21ff00",
		16#0381# => X"d4011804",
		16#0382# => X"d4012008",
		16#0383# => X"b4600010",
		16#0384# => X"00001df4",
		16#0385# => X"b4800020",
		16#0386# => X"00000000",
		16#0387# => X"00000000",
		16#0388# => X"00000000",
		16#0389# => X"00000000",
		16#038a# => X"00000000",
		16#038b# => X"00000000",
		16#038c# => X"00000000",
		16#038d# => X"00000000",
		16#038e# => X"00000000",
		16#038f# => X"00000000",
		16#0390# => X"00000000",
		16#0391# => X"00000000",
		16#0392# => X"00000000",
		16#0393# => X"00000000",
		16#0394# => X"00000000",
		16#0395# => X"00000000",
		16#0396# => X"00000000",
		16#0397# => X"00000000",
		16#0398# => X"00000000",
		16#0399# => X"00000000",
		16#039a# => X"00000000",
		16#039b# => X"00000000",
		16#039c# => X"00000000",
		16#039d# => X"00000000",
		16#039e# => X"00000000",
		16#039f# => X"00000000",
		16#03a0# => X"00000000",
		16#03a1# => X"00000000",
		16#03a2# => X"00000000",
		16#03a3# => X"00000000",
		16#03a4# => X"00000000",
		16#03a5# => X"00000000",
		16#03a6# => X"00000000",
		16#03a7# => X"00000000",
		16#03a8# => X"00000000",
		16#03a9# => X"00000000",
		16#03aa# => X"00000000",
		16#03ab# => X"00000000",
		16#03ac# => X"00000000",
		16#03ad# => X"00000000",
		16#03ae# => X"00000000",
		16#03af# => X"00000000",
		16#03b0# => X"00000000",
		16#03b1# => X"00000000",
		16#03b2# => X"00000000",
		16#03b3# => X"00000000",
		16#03b4# => X"00000000",
		16#03b5# => X"00000000",
		16#03b6# => X"00000000",
		16#03b7# => X"00000000",
		16#03b8# => X"00000000",
		16#03b9# => X"00000000",
		16#03ba# => X"00000000",
		16#03bb# => X"00000000",
		16#03bc# => X"00000000",
		16#03bd# => X"00000000",
		16#03be# => X"00000000",
		16#03bf# => X"00000000",
		16#03c0# => X"9c21ff00",
		16#03c1# => X"d4011804",
		16#03c2# => X"d4012008",
		16#03c3# => X"b4600010",
		16#03c4# => X"00001db4",
		16#03c5# => X"b4800020",
		16#03c6# => X"00000000",
		16#03c7# => X"00000000",
		16#03c8# => X"00000000",
		16#03c9# => X"00000000",
		16#03ca# => X"00000000",
		16#03cb# => X"00000000",
		16#03cc# => X"00000000",
		16#03cd# => X"00000000",
		16#03ce# => X"00000000",
		16#03cf# => X"00000000",
		16#03d0# => X"00000000",
		16#03d1# => X"00000000",
		16#03d2# => X"00000000",
		16#03d3# => X"00000000",
		16#03d4# => X"00000000",
		16#03d5# => X"00000000",
		16#03d6# => X"00000000",
		16#03d7# => X"00000000",
		16#03d8# => X"00000000",
		16#03d9# => X"00000000",
		16#03da# => X"00000000",
		16#03db# => X"00000000",
		16#03dc# => X"00000000",
		16#03dd# => X"00000000",
		16#03de# => X"00000000",
		16#03df# => X"00000000",
		16#03e0# => X"00000000",
		16#03e1# => X"00000000",
		16#03e2# => X"00000000",
		16#03e3# => X"00000000",
		16#03e4# => X"00000000",
		16#03e5# => X"00000000",
		16#03e6# => X"00000000",
		16#03e7# => X"00000000",
		16#03e8# => X"00000000",
		16#03e9# => X"00000000",
		16#03ea# => X"00000000",
		16#03eb# => X"00000000",
		16#03ec# => X"00000000",
		16#03ed# => X"00000000",
		16#03ee# => X"00000000",
		16#03ef# => X"00000000",
		16#03f0# => X"00000000",
		16#03f1# => X"00000000",
		16#03f2# => X"00000000",
		16#03f3# => X"00000000",
		16#03f4# => X"00000000",
		16#03f5# => X"00000000",
		16#03f6# => X"00000000",
		16#03f7# => X"00000000",
		16#03f8# => X"00000000",
		16#03f9# => X"00000000",
		16#03fa# => X"00000000",
		16#03fb# => X"00000000",
		16#03fc# => X"00000000",
		16#03fd# => X"00000000",
		16#03fe# => X"00000000",
		16#03ff# => X"00000000",
		16#0400# => X"9c21ff00",
		16#0401# => X"d4011804",
		16#0402# => X"d4012008",
		16#0403# => X"b4600010",
		16#0404# => X"00001d74",
		16#0405# => X"b4800020",
		16#0406# => X"00000000",
		16#0407# => X"00000000",
		16#0408# => X"00000000",
		16#0409# => X"00000000",
		16#040a# => X"00000000",
		16#040b# => X"00000000",
		16#040c# => X"00000000",
		16#040d# => X"00000000",
		16#040e# => X"00000000",
		16#040f# => X"00000000",
		16#0410# => X"00000000",
		16#0411# => X"00000000",
		16#0412# => X"00000000",
		16#0413# => X"00000000",
		16#0414# => X"00000000",
		16#0415# => X"00000000",
		16#0416# => X"00000000",
		16#0417# => X"00000000",
		16#0418# => X"00000000",
		16#0419# => X"00000000",
		16#041a# => X"00000000",
		16#041b# => X"00000000",
		16#041c# => X"00000000",
		16#041d# => X"00000000",
		16#041e# => X"00000000",
		16#041f# => X"00000000",
		16#0420# => X"00000000",
		16#0421# => X"00000000",
		16#0422# => X"00000000",
		16#0423# => X"00000000",
		16#0424# => X"00000000",
		16#0425# => X"00000000",
		16#0426# => X"00000000",
		16#0427# => X"00000000",
		16#0428# => X"00000000",
		16#0429# => X"00000000",
		16#042a# => X"00000000",
		16#042b# => X"00000000",
		16#042c# => X"00000000",
		16#042d# => X"00000000",
		16#042e# => X"00000000",
		16#042f# => X"00000000",
		16#0430# => X"00000000",
		16#0431# => X"00000000",
		16#0432# => X"00000000",
		16#0433# => X"00000000",
		16#0434# => X"00000000",
		16#0435# => X"00000000",
		16#0436# => X"00000000",
		16#0437# => X"00000000",
		16#0438# => X"00000000",
		16#0439# => X"00000000",
		16#043a# => X"00000000",
		16#043b# => X"00000000",
		16#043c# => X"00000000",
		16#043d# => X"00000000",
		16#043e# => X"00000000",
		16#043f# => X"00000000",
		16#0440# => X"9c21ff00",
		16#0441# => X"d4011804",
		16#0442# => X"d4012008",
		16#0443# => X"b4600010",
		16#0444# => X"00001d34",
		16#0445# => X"b4800020",
		16#0446# => X"00000000",
		16#0447# => X"00000000",
		16#0448# => X"00000000",
		16#0449# => X"00000000",
		16#044a# => X"00000000",
		16#044b# => X"00000000",
		16#044c# => X"00000000",
		16#044d# => X"00000000",
		16#044e# => X"00000000",
		16#044f# => X"00000000",
		16#0450# => X"00000000",
		16#0451# => X"00000000",
		16#0452# => X"00000000",
		16#0453# => X"00000000",
		16#0454# => X"00000000",
		16#0455# => X"00000000",
		16#0456# => X"00000000",
		16#0457# => X"00000000",
		16#0458# => X"00000000",
		16#0459# => X"00000000",
		16#045a# => X"00000000",
		16#045b# => X"00000000",
		16#045c# => X"00000000",
		16#045d# => X"00000000",
		16#045e# => X"00000000",
		16#045f# => X"00000000",
		16#0460# => X"00000000",
		16#0461# => X"00000000",
		16#0462# => X"00000000",
		16#0463# => X"00000000",
		16#0464# => X"00000000",
		16#0465# => X"00000000",
		16#0466# => X"00000000",
		16#0467# => X"00000000",
		16#0468# => X"00000000",
		16#0469# => X"00000000",
		16#046a# => X"00000000",
		16#046b# => X"00000000",
		16#046c# => X"00000000",
		16#046d# => X"00000000",
		16#046e# => X"00000000",
		16#046f# => X"00000000",
		16#0470# => X"00000000",
		16#0471# => X"00000000",
		16#0472# => X"00000000",
		16#0473# => X"00000000",
		16#0474# => X"00000000",
		16#0475# => X"00000000",
		16#0476# => X"00000000",
		16#0477# => X"00000000",
		16#0478# => X"00000000",
		16#0479# => X"00000000",
		16#047a# => X"00000000",
		16#047b# => X"00000000",
		16#047c# => X"00000000",
		16#047d# => X"00000000",
		16#047e# => X"00000000",
		16#047f# => X"00000000",
		16#0480# => X"9c21ff00",
		16#0481# => X"d4011804",
		16#0482# => X"d4012008",
		16#0483# => X"b4600010",
		16#0484# => X"00001cf4",
		16#0485# => X"b4800020",
		16#0486# => X"00000000",
		16#0487# => X"00000000",
		16#0488# => X"00000000",
		16#0489# => X"00000000",
		16#048a# => X"00000000",
		16#048b# => X"00000000",
		16#048c# => X"00000000",
		16#048d# => X"00000000",
		16#048e# => X"00000000",
		16#048f# => X"00000000",
		16#0490# => X"00000000",
		16#0491# => X"00000000",
		16#0492# => X"00000000",
		16#0493# => X"00000000",
		16#0494# => X"00000000",
		16#0495# => X"00000000",
		16#0496# => X"00000000",
		16#0497# => X"00000000",
		16#0498# => X"00000000",
		16#0499# => X"00000000",
		16#049a# => X"00000000",
		16#049b# => X"00000000",
		16#049c# => X"00000000",
		16#049d# => X"00000000",
		16#049e# => X"00000000",
		16#049f# => X"00000000",
		16#04a0# => X"00000000",
		16#04a1# => X"00000000",
		16#04a2# => X"00000000",
		16#04a3# => X"00000000",
		16#04a4# => X"00000000",
		16#04a5# => X"00000000",
		16#04a6# => X"00000000",
		16#04a7# => X"00000000",
		16#04a8# => X"00000000",
		16#04a9# => X"00000000",
		16#04aa# => X"00000000",
		16#04ab# => X"00000000",
		16#04ac# => X"00000000",
		16#04ad# => X"00000000",
		16#04ae# => X"00000000",
		16#04af# => X"00000000",
		16#04b0# => X"00000000",
		16#04b1# => X"00000000",
		16#04b2# => X"00000000",
		16#04b3# => X"00000000",
		16#04b4# => X"00000000",
		16#04b5# => X"00000000",
		16#04b6# => X"00000000",
		16#04b7# => X"00000000",
		16#04b8# => X"00000000",
		16#04b9# => X"00000000",
		16#04ba# => X"00000000",
		16#04bb# => X"00000000",
		16#04bc# => X"00000000",
		16#04bd# => X"00000000",
		16#04be# => X"00000000",
		16#04bf# => X"00000000",
		16#04c0# => X"9c21ff00",
		16#04c1# => X"d4011804",
		16#04c2# => X"d4012008",
		16#04c3# => X"b4600010",
		16#04c4# => X"00001cb4",
		16#04c5# => X"b4800020",
		16#04c6# => X"00000000",
		16#04c7# => X"00000000",
		16#04c8# => X"00000000",
		16#04c9# => X"00000000",
		16#04ca# => X"00000000",
		16#04cb# => X"00000000",
		16#04cc# => X"00000000",
		16#04cd# => X"00000000",
		16#04ce# => X"00000000",
		16#04cf# => X"00000000",
		16#04d0# => X"00000000",
		16#04d1# => X"00000000",
		16#04d2# => X"00000000",
		16#04d3# => X"00000000",
		16#04d4# => X"00000000",
		16#04d5# => X"00000000",
		16#04d6# => X"00000000",
		16#04d7# => X"00000000",
		16#04d8# => X"00000000",
		16#04d9# => X"00000000",
		16#04da# => X"00000000",
		16#04db# => X"00000000",
		16#04dc# => X"00000000",
		16#04dd# => X"00000000",
		16#04de# => X"00000000",
		16#04df# => X"00000000",
		16#04e0# => X"00000000",
		16#04e1# => X"00000000",
		16#04e2# => X"00000000",
		16#04e3# => X"00000000",
		16#04e4# => X"00000000",
		16#04e5# => X"00000000",
		16#04e6# => X"00000000",
		16#04e7# => X"00000000",
		16#04e8# => X"00000000",
		16#04e9# => X"00000000",
		16#04ea# => X"00000000",
		16#04eb# => X"00000000",
		16#04ec# => X"00000000",
		16#04ed# => X"00000000",
		16#04ee# => X"00000000",
		16#04ef# => X"00000000",
		16#04f0# => X"00000000",
		16#04f1# => X"00000000",
		16#04f2# => X"00000000",
		16#04f3# => X"00000000",
		16#04f4# => X"00000000",
		16#04f5# => X"00000000",
		16#04f6# => X"00000000",
		16#04f7# => X"00000000",
		16#04f8# => X"00000000",
		16#04f9# => X"00000000",
		16#04fa# => X"00000000",
		16#04fb# => X"00000000",
		16#04fc# => X"00000000",
		16#04fd# => X"00000000",
		16#04fe# => X"00000000",
		16#04ff# => X"00000000",
		16#0500# => X"9c21ff00",
		16#0501# => X"d4011804",
		16#0502# => X"d4012008",
		16#0503# => X"b4600010",
		16#0504# => X"00001c74",
		16#0505# => X"b4800020",
		16#0506# => X"00000000",
		16#0507# => X"00000000",
		16#0508# => X"00000000",
		16#0509# => X"00000000",
		16#050a# => X"00000000",
		16#050b# => X"00000000",
		16#050c# => X"00000000",
		16#050d# => X"00000000",
		16#050e# => X"00000000",
		16#050f# => X"00000000",
		16#0510# => X"00000000",
		16#0511# => X"00000000",
		16#0512# => X"00000000",
		16#0513# => X"00000000",
		16#0514# => X"00000000",
		16#0515# => X"00000000",
		16#0516# => X"00000000",
		16#0517# => X"00000000",
		16#0518# => X"00000000",
		16#0519# => X"00000000",
		16#051a# => X"00000000",
		16#051b# => X"00000000",
		16#051c# => X"00000000",
		16#051d# => X"00000000",
		16#051e# => X"00000000",
		16#051f# => X"00000000",
		16#0520# => X"00000000",
		16#0521# => X"00000000",
		16#0522# => X"00000000",
		16#0523# => X"00000000",
		16#0524# => X"00000000",
		16#0525# => X"00000000",
		16#0526# => X"00000000",
		16#0527# => X"00000000",
		16#0528# => X"00000000",
		16#0529# => X"00000000",
		16#052a# => X"00000000",
		16#052b# => X"00000000",
		16#052c# => X"00000000",
		16#052d# => X"00000000",
		16#052e# => X"00000000",
		16#052f# => X"00000000",
		16#0530# => X"00000000",
		16#0531# => X"00000000",
		16#0532# => X"00000000",
		16#0533# => X"00000000",
		16#0534# => X"00000000",
		16#0535# => X"00000000",
		16#0536# => X"00000000",
		16#0537# => X"00000000",
		16#0538# => X"00000000",
		16#0539# => X"00000000",
		16#053a# => X"00000000",
		16#053b# => X"00000000",
		16#053c# => X"00000000",
		16#053d# => X"00000000",
		16#053e# => X"00000000",
		16#053f# => X"00000000",
		16#0540# => X"9c21ff00",
		16#0541# => X"d4011804",
		16#0542# => X"d4012008",
		16#0543# => X"b4600010",
		16#0544# => X"00001c34",
		16#0545# => X"b4800020",
		16#0546# => X"00000000",
		16#0547# => X"00000000",
		16#0548# => X"00000000",
		16#0549# => X"00000000",
		16#054a# => X"00000000",
		16#054b# => X"00000000",
		16#054c# => X"00000000",
		16#054d# => X"00000000",
		16#054e# => X"00000000",
		16#054f# => X"00000000",
		16#0550# => X"00000000",
		16#0551# => X"00000000",
		16#0552# => X"00000000",
		16#0553# => X"00000000",
		16#0554# => X"00000000",
		16#0555# => X"00000000",
		16#0556# => X"00000000",
		16#0557# => X"00000000",
		16#0558# => X"00000000",
		16#0559# => X"00000000",
		16#055a# => X"00000000",
		16#055b# => X"00000000",
		16#055c# => X"00000000",
		16#055d# => X"00000000",
		16#055e# => X"00000000",
		16#055f# => X"00000000",
		16#0560# => X"00000000",
		16#0561# => X"00000000",
		16#0562# => X"00000000",
		16#0563# => X"00000000",
		16#0564# => X"00000000",
		16#0565# => X"00000000",
		16#0566# => X"00000000",
		16#0567# => X"00000000",
		16#0568# => X"00000000",
		16#0569# => X"00000000",
		16#056a# => X"00000000",
		16#056b# => X"00000000",
		16#056c# => X"00000000",
		16#056d# => X"00000000",
		16#056e# => X"00000000",
		16#056f# => X"00000000",
		16#0570# => X"00000000",
		16#0571# => X"00000000",
		16#0572# => X"00000000",
		16#0573# => X"00000000",
		16#0574# => X"00000000",
		16#0575# => X"00000000",
		16#0576# => X"00000000",
		16#0577# => X"00000000",
		16#0578# => X"00000000",
		16#0579# => X"00000000",
		16#057a# => X"00000000",
		16#057b# => X"00000000",
		16#057c# => X"00000000",
		16#057d# => X"00000000",
		16#057e# => X"00000000",
		16#057f# => X"00000000",
		16#0580# => X"9c21ff00",
		16#0581# => X"d4011804",
		16#0582# => X"d4012008",
		16#0583# => X"b4600010",
		16#0584# => X"00001bf4",
		16#0585# => X"b4800020",
		16#0586# => X"00000000",
		16#0587# => X"00000000",
		16#0588# => X"00000000",
		16#0589# => X"00000000",
		16#058a# => X"00000000",
		16#058b# => X"00000000",
		16#058c# => X"00000000",
		16#058d# => X"00000000",
		16#058e# => X"00000000",
		16#058f# => X"00000000",
		16#0590# => X"00000000",
		16#0591# => X"00000000",
		16#0592# => X"00000000",
		16#0593# => X"00000000",
		16#0594# => X"00000000",
		16#0595# => X"00000000",
		16#0596# => X"00000000",
		16#0597# => X"00000000",
		16#0598# => X"00000000",
		16#0599# => X"00000000",
		16#059a# => X"00000000",
		16#059b# => X"00000000",
		16#059c# => X"00000000",
		16#059d# => X"00000000",
		16#059e# => X"00000000",
		16#059f# => X"00000000",
		16#05a0# => X"00000000",
		16#05a1# => X"00000000",
		16#05a2# => X"00000000",
		16#05a3# => X"00000000",
		16#05a4# => X"00000000",
		16#05a5# => X"00000000",
		16#05a6# => X"00000000",
		16#05a7# => X"00000000",
		16#05a8# => X"00000000",
		16#05a9# => X"00000000",
		16#05aa# => X"00000000",
		16#05ab# => X"00000000",
		16#05ac# => X"00000000",
		16#05ad# => X"00000000",
		16#05ae# => X"00000000",
		16#05af# => X"00000000",
		16#05b0# => X"00000000",
		16#05b1# => X"00000000",
		16#05b2# => X"00000000",
		16#05b3# => X"00000000",
		16#05b4# => X"00000000",
		16#05b5# => X"00000000",
		16#05b6# => X"00000000",
		16#05b7# => X"00000000",
		16#05b8# => X"00000000",
		16#05b9# => X"00000000",
		16#05ba# => X"00000000",
		16#05bb# => X"00000000",
		16#05bc# => X"00000000",
		16#05bd# => X"00000000",
		16#05be# => X"00000000",
		16#05bf# => X"00000000",
		16#05c0# => X"9c21ff00",
		16#05c1# => X"d4011804",
		16#05c2# => X"d4012008",
		16#05c3# => X"b4600010",
		16#05c4# => X"00001bb4",
		16#05c5# => X"b4800020",
		16#05c6# => X"00000000",
		16#05c7# => X"00000000",
		16#05c8# => X"00000000",
		16#05c9# => X"00000000",
		16#05ca# => X"00000000",
		16#05cb# => X"00000000",
		16#05cc# => X"00000000",
		16#05cd# => X"00000000",
		16#05ce# => X"00000000",
		16#05cf# => X"00000000",
		16#05d0# => X"00000000",
		16#05d1# => X"00000000",
		16#05d2# => X"00000000",
		16#05d3# => X"00000000",
		16#05d4# => X"00000000",
		16#05d5# => X"00000000",
		16#05d6# => X"00000000",
		16#05d7# => X"00000000",
		16#05d8# => X"00000000",
		16#05d9# => X"00000000",
		16#05da# => X"00000000",
		16#05db# => X"00000000",
		16#05dc# => X"00000000",
		16#05dd# => X"00000000",
		16#05de# => X"00000000",
		16#05df# => X"00000000",
		16#05e0# => X"00000000",
		16#05e1# => X"00000000",
		16#05e2# => X"00000000",
		16#05e3# => X"00000000",
		16#05e4# => X"00000000",
		16#05e5# => X"00000000",
		16#05e6# => X"00000000",
		16#05e7# => X"00000000",
		16#05e8# => X"00000000",
		16#05e9# => X"00000000",
		16#05ea# => X"00000000",
		16#05eb# => X"00000000",
		16#05ec# => X"00000000",
		16#05ed# => X"00000000",
		16#05ee# => X"00000000",
		16#05ef# => X"00000000",
		16#05f0# => X"00000000",
		16#05f1# => X"00000000",
		16#05f2# => X"00000000",
		16#05f3# => X"00000000",
		16#05f4# => X"00000000",
		16#05f5# => X"00000000",
		16#05f6# => X"00000000",
		16#05f7# => X"00000000",
		16#05f8# => X"00000000",
		16#05f9# => X"00000000",
		16#05fa# => X"00000000",
		16#05fb# => X"00000000",
		16#05fc# => X"00000000",
		16#05fd# => X"00000000",
		16#05fe# => X"00000000",
		16#05ff# => X"00000000",
		16#0600# => X"9c21ff00",
		16#0601# => X"d4011804",
		16#0602# => X"d4012008",
		16#0603# => X"b4600010",
		16#0604# => X"00001b74",
		16#0605# => X"b4800020",
		16#0606# => X"00000000",
		16#0607# => X"00000000",
		16#0608# => X"00000000",
		16#0609# => X"00000000",
		16#060a# => X"00000000",
		16#060b# => X"00000000",
		16#060c# => X"00000000",
		16#060d# => X"00000000",
		16#060e# => X"00000000",
		16#060f# => X"00000000",
		16#0610# => X"00000000",
		16#0611# => X"00000000",
		16#0612# => X"00000000",
		16#0613# => X"00000000",
		16#0614# => X"00000000",
		16#0615# => X"00000000",
		16#0616# => X"00000000",
		16#0617# => X"00000000",
		16#0618# => X"00000000",
		16#0619# => X"00000000",
		16#061a# => X"00000000",
		16#061b# => X"00000000",
		16#061c# => X"00000000",
		16#061d# => X"00000000",
		16#061e# => X"00000000",
		16#061f# => X"00000000",
		16#0620# => X"00000000",
		16#0621# => X"00000000",
		16#0622# => X"00000000",
		16#0623# => X"00000000",
		16#0624# => X"00000000",
		16#0625# => X"00000000",
		16#0626# => X"00000000",
		16#0627# => X"00000000",
		16#0628# => X"00000000",
		16#0629# => X"00000000",
		16#062a# => X"00000000",
		16#062b# => X"00000000",
		16#062c# => X"00000000",
		16#062d# => X"00000000",
		16#062e# => X"00000000",
		16#062f# => X"00000000",
		16#0630# => X"00000000",
		16#0631# => X"00000000",
		16#0632# => X"00000000",
		16#0633# => X"00000000",
		16#0634# => X"00000000",
		16#0635# => X"00000000",
		16#0636# => X"00000000",
		16#0637# => X"00000000",
		16#0638# => X"00000000",
		16#0639# => X"00000000",
		16#063a# => X"00000000",
		16#063b# => X"00000000",
		16#063c# => X"00000000",
		16#063d# => X"00000000",
		16#063e# => X"00000000",
		16#063f# => X"00000000",
		16#0640# => X"9c21ff00",
		16#0641# => X"d4011804",
		16#0642# => X"d4012008",
		16#0643# => X"b4600010",
		16#0644# => X"00001b34",
		16#0645# => X"b4800020",
		16#0646# => X"00000000",
		16#0647# => X"00000000",
		16#0648# => X"00000000",
		16#0649# => X"00000000",
		16#064a# => X"00000000",
		16#064b# => X"00000000",
		16#064c# => X"00000000",
		16#064d# => X"00000000",
		16#064e# => X"00000000",
		16#064f# => X"00000000",
		16#0650# => X"00000000",
		16#0651# => X"00000000",
		16#0652# => X"00000000",
		16#0653# => X"00000000",
		16#0654# => X"00000000",
		16#0655# => X"00000000",
		16#0656# => X"00000000",
		16#0657# => X"00000000",
		16#0658# => X"00000000",
		16#0659# => X"00000000",
		16#065a# => X"00000000",
		16#065b# => X"00000000",
		16#065c# => X"00000000",
		16#065d# => X"00000000",
		16#065e# => X"00000000",
		16#065f# => X"00000000",
		16#0660# => X"00000000",
		16#0661# => X"00000000",
		16#0662# => X"00000000",
		16#0663# => X"00000000",
		16#0664# => X"00000000",
		16#0665# => X"00000000",
		16#0666# => X"00000000",
		16#0667# => X"00000000",
		16#0668# => X"00000000",
		16#0669# => X"00000000",
		16#066a# => X"00000000",
		16#066b# => X"00000000",
		16#066c# => X"00000000",
		16#066d# => X"00000000",
		16#066e# => X"00000000",
		16#066f# => X"00000000",
		16#0670# => X"00000000",
		16#0671# => X"00000000",
		16#0672# => X"00000000",
		16#0673# => X"00000000",
		16#0674# => X"00000000",
		16#0675# => X"00000000",
		16#0676# => X"00000000",
		16#0677# => X"00000000",
		16#0678# => X"00000000",
		16#0679# => X"00000000",
		16#067a# => X"00000000",
		16#067b# => X"00000000",
		16#067c# => X"00000000",
		16#067d# => X"00000000",
		16#067e# => X"00000000",
		16#067f# => X"00000000",
		16#0680# => X"9c21ff00",
		16#0681# => X"d4011804",
		16#0682# => X"d4012008",
		16#0683# => X"b4600010",
		16#0684# => X"00001af4",
		16#0685# => X"b4800020",
		16#0686# => X"00000000",
		16#0687# => X"00000000",
		16#0688# => X"00000000",
		16#0689# => X"00000000",
		16#068a# => X"00000000",
		16#068b# => X"00000000",
		16#068c# => X"00000000",
		16#068d# => X"00000000",
		16#068e# => X"00000000",
		16#068f# => X"00000000",
		16#0690# => X"00000000",
		16#0691# => X"00000000",
		16#0692# => X"00000000",
		16#0693# => X"00000000",
		16#0694# => X"00000000",
		16#0695# => X"00000000",
		16#0696# => X"00000000",
		16#0697# => X"00000000",
		16#0698# => X"00000000",
		16#0699# => X"00000000",
		16#069a# => X"00000000",
		16#069b# => X"00000000",
		16#069c# => X"00000000",
		16#069d# => X"00000000",
		16#069e# => X"00000000",
		16#069f# => X"00000000",
		16#06a0# => X"00000000",
		16#06a1# => X"00000000",
		16#06a2# => X"00000000",
		16#06a3# => X"00000000",
		16#06a4# => X"00000000",
		16#06a5# => X"00000000",
		16#06a6# => X"00000000",
		16#06a7# => X"00000000",
		16#06a8# => X"00000000",
		16#06a9# => X"00000000",
		16#06aa# => X"00000000",
		16#06ab# => X"00000000",
		16#06ac# => X"00000000",
		16#06ad# => X"00000000",
		16#06ae# => X"00000000",
		16#06af# => X"00000000",
		16#06b0# => X"00000000",
		16#06b1# => X"00000000",
		16#06b2# => X"00000000",
		16#06b3# => X"00000000",
		16#06b4# => X"00000000",
		16#06b5# => X"00000000",
		16#06b6# => X"00000000",
		16#06b7# => X"00000000",
		16#06b8# => X"00000000",
		16#06b9# => X"00000000",
		16#06ba# => X"00000000",
		16#06bb# => X"00000000",
		16#06bc# => X"00000000",
		16#06bd# => X"00000000",
		16#06be# => X"00000000",
		16#06bf# => X"00000000",
		16#06c0# => X"9c21ff00",
		16#06c1# => X"d4011804",
		16#06c2# => X"d4012008",
		16#06c3# => X"b4600010",
		16#06c4# => X"00001ab4",
		16#06c5# => X"b4800020",
		16#06c6# => X"00000000",
		16#06c7# => X"00000000",
		16#06c8# => X"00000000",
		16#06c9# => X"00000000",
		16#06ca# => X"00000000",
		16#06cb# => X"00000000",
		16#06cc# => X"00000000",
		16#06cd# => X"00000000",
		16#06ce# => X"00000000",
		16#06cf# => X"00000000",
		16#06d0# => X"00000000",
		16#06d1# => X"00000000",
		16#06d2# => X"00000000",
		16#06d3# => X"00000000",
		16#06d4# => X"00000000",
		16#06d5# => X"00000000",
		16#06d6# => X"00000000",
		16#06d7# => X"00000000",
		16#06d8# => X"00000000",
		16#06d9# => X"00000000",
		16#06da# => X"00000000",
		16#06db# => X"00000000",
		16#06dc# => X"00000000",
		16#06dd# => X"00000000",
		16#06de# => X"00000000",
		16#06df# => X"00000000",
		16#06e0# => X"00000000",
		16#06e1# => X"00000000",
		16#06e2# => X"00000000",
		16#06e3# => X"00000000",
		16#06e4# => X"00000000",
		16#06e5# => X"00000000",
		16#06e6# => X"00000000",
		16#06e7# => X"00000000",
		16#06e8# => X"00000000",
		16#06e9# => X"00000000",
		16#06ea# => X"00000000",
		16#06eb# => X"00000000",
		16#06ec# => X"00000000",
		16#06ed# => X"00000000",
		16#06ee# => X"00000000",
		16#06ef# => X"00000000",
		16#06f0# => X"00000000",
		16#06f1# => X"00000000",
		16#06f2# => X"00000000",
		16#06f3# => X"00000000",
		16#06f4# => X"00000000",
		16#06f5# => X"00000000",
		16#06f6# => X"00000000",
		16#06f7# => X"00000000",
		16#06f8# => X"00000000",
		16#06f9# => X"00000000",
		16#06fa# => X"00000000",
		16#06fb# => X"00000000",
		16#06fc# => X"00000000",
		16#06fd# => X"00000000",
		16#06fe# => X"00000000",
		16#06ff# => X"00000000",
		16#0700# => X"9c21ff00",
		16#0701# => X"d4011804",
		16#0702# => X"d4012008",
		16#0703# => X"b4600010",
		16#0704# => X"00001a74",
		16#0705# => X"b4800020",
		16#0706# => X"00000000",
		16#0707# => X"00000000",
		16#0708# => X"00000000",
		16#0709# => X"00000000",
		16#070a# => X"00000000",
		16#070b# => X"00000000",
		16#070c# => X"00000000",
		16#070d# => X"00000000",
		16#070e# => X"00000000",
		16#070f# => X"00000000",
		16#0710# => X"00000000",
		16#0711# => X"00000000",
		16#0712# => X"00000000",
		16#0713# => X"00000000",
		16#0714# => X"00000000",
		16#0715# => X"00000000",
		16#0716# => X"00000000",
		16#0717# => X"00000000",
		16#0718# => X"00000000",
		16#0719# => X"00000000",
		16#071a# => X"00000000",
		16#071b# => X"00000000",
		16#071c# => X"00000000",
		16#071d# => X"00000000",
		16#071e# => X"00000000",
		16#071f# => X"00000000",
		16#0720# => X"00000000",
		16#0721# => X"00000000",
		16#0722# => X"00000000",
		16#0723# => X"00000000",
		16#0724# => X"00000000",
		16#0725# => X"00000000",
		16#0726# => X"00000000",
		16#0727# => X"00000000",
		16#0728# => X"00000000",
		16#0729# => X"00000000",
		16#072a# => X"00000000",
		16#072b# => X"00000000",
		16#072c# => X"00000000",
		16#072d# => X"00000000",
		16#072e# => X"00000000",
		16#072f# => X"00000000",
		16#0730# => X"00000000",
		16#0731# => X"00000000",
		16#0732# => X"00000000",
		16#0733# => X"00000000",
		16#0734# => X"00000000",
		16#0735# => X"00000000",
		16#0736# => X"00000000",
		16#0737# => X"00000000",
		16#0738# => X"00000000",
		16#0739# => X"00000000",
		16#073a# => X"00000000",
		16#073b# => X"00000000",
		16#073c# => X"00000000",
		16#073d# => X"00000000",
		16#073e# => X"00000000",
		16#073f# => X"00000000",
		16#0740# => X"9c21ff00",
		16#0741# => X"d4011804",
		16#0742# => X"d4012008",
		16#0743# => X"b4600010",
		16#0744# => X"00001a34",
		16#0745# => X"b4800020",
		16#0746# => X"00000000",
		16#0747# => X"00000000",
		16#0748# => X"00000000",
		16#0749# => X"00000000",
		16#074a# => X"00000000",
		16#074b# => X"00000000",
		16#074c# => X"00000000",
		16#074d# => X"00000000",
		16#074e# => X"00000000",
		16#074f# => X"00000000",
		16#0750# => X"00000000",
		16#0751# => X"00000000",
		16#0752# => X"00000000",
		16#0753# => X"00000000",
		16#0754# => X"00000000",
		16#0755# => X"00000000",
		16#0756# => X"00000000",
		16#0757# => X"00000000",
		16#0758# => X"00000000",
		16#0759# => X"00000000",
		16#075a# => X"00000000",
		16#075b# => X"00000000",
		16#075c# => X"00000000",
		16#075d# => X"00000000",
		16#075e# => X"00000000",
		16#075f# => X"00000000",
		16#0760# => X"00000000",
		16#0761# => X"00000000",
		16#0762# => X"00000000",
		16#0763# => X"00000000",
		16#0764# => X"00000000",
		16#0765# => X"00000000",
		16#0766# => X"00000000",
		16#0767# => X"00000000",
		16#0768# => X"00000000",
		16#0769# => X"00000000",
		16#076a# => X"00000000",
		16#076b# => X"00000000",
		16#076c# => X"00000000",
		16#076d# => X"00000000",
		16#076e# => X"00000000",
		16#076f# => X"00000000",
		16#0770# => X"00000000",
		16#0771# => X"00000000",
		16#0772# => X"00000000",
		16#0773# => X"00000000",
		16#0774# => X"00000000",
		16#0775# => X"00000000",
		16#0776# => X"00000000",
		16#0777# => X"00000000",
		16#0778# => X"00000000",
		16#0779# => X"00000000",
		16#077a# => X"00000000",
		16#077b# => X"00000000",
		16#077c# => X"00000000",
		16#077d# => X"00000000",
		16#077e# => X"00000000",
		16#077f# => X"00000000",
		16#0780# => X"9c21ff00",
		16#0781# => X"d4011804",
		16#0782# => X"d4012008",
		16#0783# => X"b4600010",
		16#0784# => X"000019f4",
		16#0785# => X"b4800020",
		16#0786# => X"00000000",
		16#0787# => X"00000000",
		16#0788# => X"00000000",
		16#0789# => X"00000000",
		16#078a# => X"00000000",
		16#078b# => X"00000000",
		16#078c# => X"00000000",
		16#078d# => X"00000000",
		16#078e# => X"00000000",
		16#078f# => X"00000000",
		16#0790# => X"00000000",
		16#0791# => X"00000000",
		16#0792# => X"00000000",
		16#0793# => X"00000000",
		16#0794# => X"00000000",
		16#0795# => X"00000000",
		16#0796# => X"00000000",
		16#0797# => X"00000000",
		16#0798# => X"00000000",
		16#0799# => X"00000000",
		16#079a# => X"00000000",
		16#079b# => X"00000000",
		16#079c# => X"00000000",
		16#079d# => X"00000000",
		16#079e# => X"00000000",
		16#079f# => X"00000000",
		16#07a0# => X"00000000",
		16#07a1# => X"00000000",
		16#07a2# => X"00000000",
		16#07a3# => X"00000000",
		16#07a4# => X"00000000",
		16#07a5# => X"00000000",
		16#07a6# => X"00000000",
		16#07a7# => X"00000000",
		16#07a8# => X"00000000",
		16#07a9# => X"00000000",
		16#07aa# => X"00000000",
		16#07ab# => X"00000000",
		16#07ac# => X"00000000",
		16#07ad# => X"00000000",
		16#07ae# => X"00000000",
		16#07af# => X"00000000",
		16#07b0# => X"00000000",
		16#07b1# => X"00000000",
		16#07b2# => X"00000000",
		16#07b3# => X"00000000",
		16#07b4# => X"00000000",
		16#07b5# => X"00000000",
		16#07b6# => X"00000000",
		16#07b7# => X"00000000",
		16#07b8# => X"00000000",
		16#07b9# => X"00000000",
		16#07ba# => X"00000000",
		16#07bb# => X"00000000",
		16#07bc# => X"00000000",
		16#07bd# => X"00000000",
		16#07be# => X"00000000",
		16#07bf# => X"00000000",
		16#07c0# => X"9c21ff00",
		16#07c1# => X"d4011804",
		16#07c2# => X"d4012008",
		16#07c3# => X"b4600010",
		16#07c4# => X"000019b4",
		16#07c5# => X"b4800020",
		16#07c6# => X"00000000",
		16#07c7# => X"00000000",
		16#07c8# => X"00000000",
		16#07c9# => X"00000000",
		16#07ca# => X"00000000",
		16#07cb# => X"00000000",
		16#07cc# => X"00000000",
		16#07cd# => X"00000000",
		16#07ce# => X"00000000",
		16#07cf# => X"00000000",
		16#07d0# => X"00000000",
		16#07d1# => X"00000000",
		16#07d2# => X"00000000",
		16#07d3# => X"00000000",
		16#07d4# => X"00000000",
		16#07d5# => X"00000000",
		16#07d6# => X"00000000",
		16#07d7# => X"00000000",
		16#07d8# => X"00000000",
		16#07d9# => X"00000000",
		16#07da# => X"00000000",
		16#07db# => X"00000000",
		16#07dc# => X"00000000",
		16#07dd# => X"00000000",
		16#07de# => X"00000000",
		16#07df# => X"00000000",
		16#07e0# => X"00000000",
		16#07e1# => X"00000000",
		16#07e2# => X"00000000",
		16#07e3# => X"00000000",
		16#07e4# => X"00000000",
		16#07e5# => X"00000000",
		16#07e6# => X"00000000",
		16#07e7# => X"00000000",
		16#07e8# => X"00000000",
		16#07e9# => X"00000000",
		16#07ea# => X"00000000",
		16#07eb# => X"00000000",
		16#07ec# => X"00000000",
		16#07ed# => X"00000000",
		16#07ee# => X"00000000",
		16#07ef# => X"00000000",
		16#07f0# => X"00000000",
		16#07f1# => X"00000000",
		16#07f2# => X"00000000",
		16#07f3# => X"00000000",
		16#07f4# => X"00000000",
		16#07f5# => X"00000000",
		16#07f6# => X"00000000",
		16#07f7# => X"00000000",
		16#07f8# => X"00000000",
		16#07f9# => X"00000000",
		16#07fa# => X"00000000",
		16#07fb# => X"00000000",
		16#07fc# => X"00000000",
		16#07fd# => X"00000000",
		16#07fe# => X"00000000",
		16#07ff# => X"15000000",
		16#0800# => X"15000000",
		16#0801# => X"9c21fffc",
		16#0802# => X"d4014800",
		16#0803# => X"04000071",
		16#0804# => X"15000000",
		16#0805# => X"04004660",
		16#0806# => X"15000000",
		16#0807# => X"85210000",
		16#0808# => X"44004800",
		16#0809# => X"9c210004",
		16#080a# => X"18200001",
		16#080b# => X"a82138f0",
		16#080c# => X"84210000",
		16#080d# => X"18400001",
		16#080e# => X"a84238f4",
		16#080f# => X"84420000",
		16#0810# => X"e0211000",
		16#0811# => X"e0410804",
		16#0812# => X"b460c002",
		16#0813# => X"b0838000",
		16#0814# => X"e0212000",
		16#0815# => X"18600001",
		16#0816# => X"a86363d8",
		16#0817# => X"d4030800",
		16#0818# => X"040018b2",
		16#0819# => X"15000000",
		16#081a# => X"18600001",
		16#081b# => X"a8636ddc",
		16#081c# => X"18800001",
		16#081d# => X"a8849ad4",
		16#081e# => X"d4030000",
		16#081f# => X"e4832000",
		16#0820# => X"13fffffe",
		16#0821# => X"9c630004",
		16#0822# => X"0400449b",
		16#0823# => X"15000000",
		16#0824# => X"07ffffdd",
		16#0825# => X"15000000",
		16#0826# => X"18600001",
		16#0827# => X"04001605",
		16#0828# => X"a86339f8",
		16#0829# => X"18800001",
		16#082a# => X"a88438fc",
		16#082b# => X"84840000",
		16#082c# => X"e4240000",
		16#082d# => X"0c000004",
		16#082e# => X"e0600004",
		16#082f# => X"04004586",
		16#0830# => X"15000000",
		16#0831# => X"e0600004",
		16#0832# => X"e0800004",
		16#0833# => X"04000084",
		16#0834# => X"e0a00004",
		16#0835# => X"04001600",
		16#0836# => X"9c6b0000",
		16#0837# => X"00000000",
		16#0838# => X"15000000",
		16#0839# => X"d7e187f8",
		16#083a# => X"1a000001",
		16#083b# => X"d7e117f0",
		16#083c# => X"aa106ddc",
		16#083d# => X"d7e14ffc",
		16#083e# => X"8c500000",
		16#083f# => X"d7e177f4",
		16#0840# => X"bc220000",
		16#0841# => X"10000027",
		16#0842# => X"9c21fff0",
		16#0843# => X"19c00001",
		16#0844# => X"18800001",
		16#0845# => X"a9ce63d0",
		16#0846# => X"a88463cc",
		16#0847# => X"18400001",
		16#0848# => X"e1ce2002",
		16#0849# => X"a8426de0",
		16#084a# => X"b9ce0082",
		16#084b# => X"84620000",
		16#084c# => X"9dceffff",
		16#084d# => X"e4637000",
		16#084e# => X"10000010",
		16#084f# => X"15000000",
		16#0850# => X"9c630001",
		16#0851# => X"18a00001",
		16#0852# => X"b8830002",
		16#0853# => X"a8a563cc",
		16#0854# => X"d4021800",
		16#0855# => X"e0642800",
		16#0856# => X"84630000",
		16#0857# => X"48001800",
		16#0858# => X"15000000",
		16#0859# => X"84620000",
		16#085a# => X"e4837000",
		16#085b# => X"13fffff6",
		16#085c# => X"9c630001",
		16#085d# => X"9c63ffff",
		16#085e# => X"18400000",
		16#085f# => X"a8420000",
		16#0860# => X"bc020000",
		16#0861# => X"10000006",
		16#0862# => X"9c400001",
		16#0863# => X"18600001",
		16#0864# => X"07fff79c",
		16#0865# => X"a86343c0",
		16#0866# => X"9c400001",
		16#0867# => X"d8101000",
		16#0868# => X"9c210010",
		16#0869# => X"8521fffc",
		16#086a# => X"8441fff0",
		16#086b# => X"85c1fff4",
		16#086c# => X"44004800",
		16#086d# => X"8601fff8",
		16#086e# => X"d7e14ffc",
		16#086f# => X"9c21fffc",
		16#0870# => X"9c210004",
		16#0871# => X"8521fffc",
		16#0872# => X"44004800",
		16#0873# => X"15000000",
		16#0874# => X"18600000",
		16#0875# => X"d7e14ffc",
		16#0876# => X"a8630000",
		16#0877# => X"bc030000",
		16#0878# => X"10000007",
		16#0879# => X"9c21fffc",
		16#087a# => X"18600001",
		16#087b# => X"18800001",
		16#087c# => X"a86343c0",
		16#087d# => X"07fff783",
		16#087e# => X"a8846de4",
		16#087f# => X"18600001",
		16#0880# => X"a86363d4",
		16#0881# => X"84830000",
		16#0882# => X"bc040000",
		16#0883# => X"1000000a",
		16#0884# => X"18800000",
		16#0885# => X"a8840000",
		16#0886# => X"bc040000",
		16#0887# => X"10000006",
		16#0888# => X"15000000",
		16#0889# => X"9c210004",
		16#088a# => X"8521fffc",
		16#088b# => X"44002000",
		16#088c# => X"15000000",
		16#088d# => X"9c210004",
		16#088e# => X"8521fffc",
		16#088f# => X"44004800",
		16#0890# => X"15000000",
		16#0891# => X"d7e14ffc",
		16#0892# => X"9c21fffc",
		16#0893# => X"9c210004",
		16#0894# => X"8521fffc",
		16#0895# => X"44004800",
		16#0896# => X"15000000",
		16#0897# => X"85630000",
		16#0898# => X"84640000",
		16#0899# => X"44004800",
		16#089a# => X"e16b1802",
		16#089b# => X"9d600001",
		16#089c# => X"d7e117fc",
		16#089d# => X"e0a35800",
		16#089e# => X"e0841802",
		16#089f# => X"e4652000",
		16#08a0# => X"10000014",
		16#08a1# => X"9c21fffc",
		16#08a2# => X"18400001",
		16#08a3# => X"b8c30002",
		16#08a4# => X"a8428ac8",
		16#08a5# => X"b8650002",
		16#08a6# => X"e0c61000",
		16#08a7# => X"e0631000",
		16#08a8# => X"85060000",
		16#08a9# => X"84c30000",
		16#08aa# => X"9ca50001",
		16#08ab# => X"e5483000",
		16#08ac# => X"10000003",
		16#08ad# => X"9ce00000",
		16#08ae# => X"a8eb0000",
		16#08af# => X"9c630004",
		16#08b0# => X"a9670000",
		16#08b1# => X"e4852000",
		16#08b2# => X"13fffff7",
		16#08b3# => X"a9060000",
		16#08b4# => X"9c210004",
		16#08b5# => X"44004800",
		16#08b6# => X"8441fffc",
		16#08b7# => X"d7e14ffc",
		16#08b8# => X"d7e197e4",
		16#08b9# => X"d7e1c7f0",
		16#08ba# => X"d7e117d8",
		16#08bb# => X"d7e177dc",
		16#08bc# => X"d7e187e0",
		16#08bd# => X"d7e1a7e8",
		16#08be# => X"d7e1b7ec",
		16#08bf# => X"d7e1d7f4",
		16#08c0# => X"d7e1e7f8",
		16#08c1# => X"04000153",
		16#08c2# => X"9c21ffd4",
		16#08c3# => X"04000157",
		16#08c4# => X"aa4b0000",
		16#08c5# => X"bc2b0000",
		16#08c6# => X"0c000078",
		16#08c7# => X"ab0b0000",
		16#08c8# => X"1a800001",
		16#08c9# => X"9c600000",
		16#08ca# => X"04000156",
		16#08cb# => X"aa948ac4",
		16#08cc# => X"b878000a",
		16#08cd# => X"04000a33",
		16#08ce# => X"a8920000",
		16#08cf# => X"18a00001",
		16#08d0# => X"b96b0002",
		16#08d1# => X"a8a58ac8",
		16#08d2# => X"9c600400",
		16#08d3# => X"a8920000",
		16#08d4# => X"04000a2c",
		16#08d5# => X"e04b2800",
		16#08d6# => X"18c00000",
		16#08d7# => X"a8620000",
		16#08d8# => X"a88b0000",
		16#08d9# => X"9ca00004",
		16#08da# => X"a8c6225c",
		16#08db# => X"040019c0",
		16#08dc# => X"9c52ffff",
		16#08dd# => X"e5781000",
		16#08de# => X"0c00005c",
		16#08df# => X"15000000",
		16#08e0# => X"bc380000",
		16#08e1# => X"10000047",
		16#08e2# => X"1860f000",
		16#08e3# => X"a8980000",
		16#08e4# => X"040000ed",
		16#08e5# => X"1b800001",
		16#08e6# => X"18600001",
		16#08e7# => X"ab9c8abc",
		16#08e8# => X"a8633a99",
		16#08e9# => X"04001965",
		16#08ea# => X"d41c5800",
		16#08eb# => X"bdb20000",
		16#08ec# => X"10000028",
		16#08ed# => X"bb52000a",
		16#08ee# => X"86d40000",
		16#08ef# => X"a9d80000",
		16#08f0# => X"a86e0000",
		16#08f1# => X"a8920000",
		16#08f2# => X"04000a0e",
		16#08f3# => X"9dce0400",
		16#08f4# => X"a86e0000",
		16#08f5# => X"aa0b0000",
		16#08f6# => X"a8920000",
		16#08f7# => X"04000a09",
		16#08f8# => X"9c4b0001",
		16#08f9# => X"e16b8002",
		16#08fa# => X"9dabffff",
		16#08fb# => X"e4626800",
		16#08fc# => X"10000014",
		16#08fd# => X"9ce00001",
		16#08fe# => X"18800001",
		16#08ff# => X"b8700002",
		16#0900# => X"a8848ac8",
		16#0901# => X"b8a20002",
		16#0902# => X"e0632000",
		16#0903# => X"e0a52000",
		16#0904# => X"85030000",
		16#0905# => X"85850000",
		16#0906# => X"9c420001",
		16#0907# => X"e5486000",
		16#0908# => X"9cc00000",
		16#0909# => X"10000003",
		16#090a# => X"a90c0000",
		16#090b# => X"a8c70000",
		16#090c# => X"9ca50004",
		16#090d# => X"e4826800",
		16#090e# => X"13fffff7",
		16#090f# => X"a8e60000",
		16#0910# => X"e42ed000",
		16#0911# => X"13ffffdf",
		16#0912# => X"e2d63800",
		16#0913# => X"d414b000",
		16#0914# => X"84540000",
		16#0915# => X"e4229000",
		16#0916# => X"0c000080",
		16#0917# => X"15000000",
		16#0918# => X"18600001",
		16#0919# => X"04001978",
		16#091a# => X"a8633aca",
		16#091b# => X"18400001",
		16#091c# => X"849c0000",
		16#091d# => X"a8428ac0",
		16#091e# => X"18600001",
		16#091f# => X"84420000",
		16#0920# => X"a8633af4",
		16#0921# => X"e0441002",
		16#0922# => X"0400192c",
		16#0923# => X"d4011000",
		16#0924# => X"04000107",
		16#0925# => X"9c600000",
		16#0926# => X"00000007",
		16#0927# => X"9c21002c",
		16#0928# => X"04000103",
		16#0929# => X"a8780000",
		16#092a# => X"040000f6",
		16#092b# => X"9c600000",
		16#092c# => X"9c21002c",
		16#092d# => X"85740000",
		16#092e# => X"8521fffc",
		16#092f# => X"9d6bffff",
		16#0930# => X"8441ffd8",
		16#0931# => X"85c1ffdc",
		16#0932# => X"8601ffe0",
		16#0933# => X"8641ffe4",
		16#0934# => X"8681ffe8",
		16#0935# => X"86c1ffec",
		16#0936# => X"8701fff0",
		16#0937# => X"8741fff4",
		16#0938# => X"44004800",
		16#0939# => X"8781fff8",
		16#093a# => X"040000e6",
		16#093b# => X"9c780001",
		16#093c# => X"03ffffa5",
		16#093d# => X"bc380000",
		16#093e# => X"1860017d",
		16#093f# => X"1a800001",
		16#0940# => X"a8637840",
		16#0941# => X"0400005a",
		16#0942# => X"9c400001",
		16#0943# => X"18600001",
		16#0944# => X"9c800400",
		16#0945# => X"a8633a14",
		16#0946# => X"aa948ac4",
		16#0947# => X"d4012000",
		16#0948# => X"04001906",
		16#0949# => X"d4141000",
		16#094a# => X"04001bda",
		16#094b# => X"15000000",
		16#094c# => X"bc6bffff",
		16#094d# => X"0c000047",
		16#094e# => X"15000000",
		16#094f# => X"18600001",
		16#0950# => X"e04b1000",
		16#0951# => X"a8638ac8",
		16#0952# => X"9e000000",
		16#0953# => X"19c00001",
		16#0954# => X"9e100001",
		16#0955# => X"d4031000",
		16#0956# => X"bc300400",
		16#0957# => X"0c000015",
		16#0958# => X"a9ce8acc",
		16#0959# => X"04001bcb",
		16#095a# => X"9c400001",
		16#095b# => X"bc6bffff",
		16#095c# => X"10000004",
		16#095d# => X"e04b1000",
		16#095e# => X"9c400000",
		16#095f# => X"e04b1000",
		16#0960# => X"bc100001",
		16#0961# => X"10000007",
		16#0962# => X"d40e1000",
		16#0963# => X"84aefffc",
		16#0964# => X"e5622800",
		16#0965# => X"10000003",
		16#0966# => X"9c400000",
		16#0967# => X"d4141000",
		16#0968# => X"9e100001",
		16#0969# => X"bc300400",
		16#096a# => X"13ffffef",
		16#096b# => X"9dce0004",
		16#096c# => X"84540000",
		16#096d# => X"bc020000",
		16#096e# => X"0c000021",
		16#096f# => X"15000000",
		16#0970# => X"18600001",
		16#0971# => X"04001920",
		16#0972# => X"a8633a5c",
		16#0973# => X"18600001",
		16#0974# => X"d4019000",
		16#0975# => X"a8633a74",
		16#0976# => X"040018d8",
		16#0977# => X"18400001",
		16#0978# => X"1860f000",
		16#0979# => X"9c800000",
		16#097a# => X"04000025",
		16#097b# => X"a8428ac0",
		16#097c# => X"1860f000",
		16#097d# => X"04000028",
		16#097e# => X"9c800000",
		16#097f# => X"9ca00002",
		16#0980# => X"1860f000",
		16#0981# => X"04000038",
		16#0982# => X"9c800000",
		16#0983# => X"9c800000",
		16#0984# => X"0400004d",
		16#0985# => X"1860f000",
		16#0986# => X"9c600000",
		16#0987# => X"040000a4",
		16#0988# => X"d4025800",
		16#0989# => X"04000097",
		16#098a# => X"9c600000",
		16#098b# => X"040000a9",
		16#098c# => X"9c600000",
		16#098d# => X"03ffff40",
		16#098e# => X"b878000a",
		16#098f# => X"18600001",
		16#0990# => X"04001901",
		16#0991# => X"a8633a3c",
		16#0992# => X"03ffffe2",
		16#0993# => X"18600001",
		16#0994# => X"03ffffbb",
		16#0995# => X"a8580000",
		16#0996# => X"18600001",
		16#0997# => X"040018fa",
		16#0998# => X"a8633aad",
		16#0999# => X"03ffff83",
		16#099a# => X"18400001",
		16#099b# => X"18800001",
		16#099c# => X"a8846e7c",
		16#099d# => X"44004800",
		16#099e# => X"d4041800",
		16#099f# => X"b8840004",
		16#09a0# => X"e0641800",
		16#09a1# => X"9c800001",
		16#09a2# => X"d4032000",
		16#09a3# => X"44004800",
		16#09a4# => X"15000000",
		16#09a5# => X"b8840004",
		16#09a6# => X"e0641800",
		16#09a7# => X"9c800002",
		16#09a8# => X"d4032000",
		16#09a9# => X"44004800",
		16#09aa# => X"15000000",
		16#09ab# => X"b8840004",
		16#09ac# => X"d7e117fc",
		16#09ad# => X"9c400000",
		16#09ae# => X"e0641800",
		16#09af# => X"9c21fffc",
		16#09b0# => X"d4031000",
		16#09b1# => X"9c210004",
		16#09b2# => X"44004800",
		16#09b3# => X"8441fffc",
		16#09b4# => X"b8840004",
		16#09b5# => X"e0632000",
		16#09b6# => X"85630004",
		16#09b7# => X"44004800",
		16#09b8# => X"15000000",
		16#09b9# => X"b8c40004",
		16#09ba# => X"9c630004",
		16#09bb# => X"d7e117fc",
		16#09bc# => X"e0633000",
		16#09bd# => X"9c21fffc",
		16#09be# => X"d4032800",
		16#09bf# => X"9d60ffff",
		16#09c0# => X"84630000",
		16#09c1# => X"e4232800",
		16#09c2# => X"10000007",
		16#09c3# => X"b8840002",
		16#09c4# => X"18400001",
		16#09c5# => X"a8426dfc",
		16#09c6# => X"9d600000",
		16#09c7# => X"e0841000",
		16#09c8# => X"d4041800",
		16#09c9# => X"9c210004",
		16#09ca# => X"44004800",
		16#09cb# => X"8441fffc",
		16#09cc# => X"b8840004",
		16#09cd# => X"e0632000",
		16#09ce# => X"85630008",
		16#09cf# => X"44004800",
		16#09d0# => X"15000000",
		16#09d1# => X"18a00001",
		16#09d2# => X"d7e117f4",
		16#09d3# => X"b8440002",
		16#09d4# => X"a8a56dfc",
		16#09d5# => X"d7e14ffc",
		16#09d6# => X"e0422800",
		16#09d7# => X"d7e177f8",
		16#09d8# => X"84420000",
		16#09d9# => X"bc020000",
		16#09da# => X"0c000003",
		16#09db# => X"9c21fff4",
		16#09dc# => X"9c400001",
		16#09dd# => X"b8a40004",
		16#09de# => X"9c8003e8",
		16#09df# => X"e0a32800",
		16#09e0# => X"18600001",
		16#09e1# => X"85c50008",
		16#09e2# => X"a8636e7c",
		16#09e3# => X"0400091d",
		16#09e4# => X"84630000",
		16#09e5# => X"a86e0000",
		16#09e6# => X"040008db",
		16#09e7# => X"a88b0000",
		16#09e8# => X"9c21000c",
		16#09e9# => X"e1625b06",
		16#09ea# => X"8521fffc",
		16#09eb# => X"8441fff4",
		16#09ec# => X"44004800",
		16#09ed# => X"85c1fff8",
		16#09ee# => X"b8840004",
		16#09ef# => X"e0632000",
		16#09f0# => X"84630008",
		16#09f1# => X"44004800",
		16#09f2# => X"d4051800",
		16#09f3# => X"d7e177f4",
		16#09f4# => X"a9c50000",
		16#09f5# => X"18a00001",
		16#09f6# => X"d7e117f0",
		16#09f7# => X"b8440002",
		16#09f8# => X"a8a56dfc",
		16#09f9# => X"d7e14ffc",
		16#09fa# => X"e0422800",
		16#09fb# => X"d7e187f8",
		16#09fc# => X"84420000",
		16#09fd# => X"bc020000",
		16#09fe# => X"0c000003",
		16#09ff# => X"9c21fff0",
		16#0a00# => X"9c400001",
		16#0a01# => X"b8a40004",
		16#0a02# => X"9c8003e8",
		16#0a03# => X"e0a32800",
		16#0a04# => X"18600001",
		16#0a05# => X"86050008",
		16#0a06# => X"a8636e7c",
		16#0a07# => X"040008f9",
		16#0a08# => X"84630000",
		16#0a09# => X"a8700000",
		16#0a0a# => X"040008b7",
		16#0a0b# => X"a88b0000",
		16#0a0c# => X"e0425b06",
		16#0a0d# => X"d40e1000",
		16#0a0e# => X"9c210010",
		16#0a0f# => X"8521fffc",
		16#0a10# => X"8441fff0",
		16#0a11# => X"85c1fff4",
		16#0a12# => X"44004800",
		16#0a13# => X"8601fff8",
		16#0a14# => X"d7e14ffc",
		16#0a15# => X"9c21fffc",
		16#0a16# => X"9c210004",
		16#0a17# => X"8521fffc",
		16#0a18# => X"000017d3",
		16#0a19# => X"a860c000",
		16#0a1a# => X"d7e14ffc",
		16#0a1b# => X"9c21fffc",
		16#0a1c# => X"9c210004",
		16#0a1d# => X"8521fffc",
		16#0a1e# => X"000017cd",
		16#0a1f# => X"a860c002",
		16#0a20# => X"9c800001",
		16#0a21# => X"18a00001",
		16#0a22# => X"e0641808",
		16#0a23# => X"a8a56e80",
		16#0a24# => X"84850000",
		16#0a25# => X"e0832003",
		16#0a26# => X"bc040000",
		16#0a27# => X"13fffffd",
		16#0a28# => X"15000000",
		16#0a29# => X"44004800",
		16#0a2a# => X"15000000",
		16#0a2b# => X"18800001",
		16#0a2c# => X"9ca00001",
		16#0a2d# => X"a8846e80",
		16#0a2e# => X"e0651808",
		16#0a2f# => X"84a40000",
		16#0a30# => X"e0632804",
		16#0a31# => X"d4041800",
		16#0a32# => X"44004800",
		16#0a33# => X"15000000",
		16#0a34# => X"9ca00001",
		16#0a35# => X"18800001",
		16#0a36# => X"e0651808",
		16#0a37# => X"a8846e80",
		16#0a38# => X"ac63ffff",
		16#0a39# => X"84a40000",
		16#0a3a# => X"e0632803",
		16#0a3b# => X"d4041800",
		16#0a3c# => X"44004800",
		16#0a3d# => X"15000000",
		16#0a3e# => X"18600001",
		16#0a3f# => X"d7e117fc",
		16#0a40# => X"a8636e80",
		16#0a41# => X"9c400000",
		16#0a42# => X"9c21fffc",
		16#0a43# => X"d4031000",
		16#0a44# => X"9c210004",
		16#0a45# => X"44004800",
		16#0a46# => X"8441fffc",
		16#0a47# => X"18600001",
		16#0a48# => X"9c80ffff",
		16#0a49# => X"a8636e80",
		16#0a4a# => X"d4032000",
		16#0a4b# => X"44004800",
		16#0a4c# => X"15000000",
		16#0a4d# => X"d7e14ffc",
		16#0a4e# => X"9c21fffc",
		16#0a4f# => X"a860c800",
		16#0a50# => X"9c210004",
		16#0a51# => X"8521fffc",
		16#0a52# => X"00001796",
		16#0a53# => X"9c800001",
		16#0a54# => X"d7e14ffc",
		16#0a55# => X"9c21fffc",
		16#0a56# => X"a860c800",
		16#0a57# => X"9c210004",
		16#0a58# => X"8521fffc",
		16#0a59# => X"0000178f",
		16#0a5a# => X"9c800000",
		16#0a5b# => X"d7e177f8",
		16#0a5c# => X"a9c40000",
		16#0a5d# => X"a880c83e",
		16#0a5e# => X"d7e14ffc",
		16#0a5f# => X"d7e117f4",
		16#0a60# => X"9c21fff4",
		16#0a61# => X"a8430000",
		16#0a62# => X"04001789",
		16#0a63# => X"e06e2000",
		16#0a64# => X"a880c83c",
		16#0a65# => X"d4025800",
		16#0a66# => X"04001785",
		16#0a67# => X"e06e2000",
		16#0a68# => X"a880c83d",
		16#0a69# => X"9d6b0001",
		16#0a6a# => X"e06e2000",
		16#0a6b# => X"04001780",
		16#0a6c# => X"d4025804",
		16#0a6d# => X"a880c83f",
		16#0a6e# => X"9d6b0001",
		16#0a6f# => X"e06e2000",
		16#0a70# => X"0400177b",
		16#0a71# => X"d402580c",
		16#0a72# => X"a86b0000",
		16#0a73# => X"04000c58",
		16#0a74# => X"d4025810",
		16#0a75# => X"84620000",
		16#0a76# => X"04000c55",
		16#0a77# => X"a9cb0000",
		16#0a78# => X"a86e0000",
		16#0a79# => X"04000aa7",
		16#0a7a# => X"a88b0000",
		16#0a7b# => X"d4025808",
		16#0a7c# => X"9c21000c",
		16#0a7d# => X"8521fffc",
		16#0a7e# => X"8441fff4",
		16#0a7f# => X"44004800",
		16#0a80# => X"85c1fff8",
		16#0a81# => X"d7e14ffc",
		16#0a82# => X"d7e117d4",
		16#0a83# => X"d7e177d8",
		16#0a84# => X"d7e187dc",
		16#0a85# => X"d7e197e0",
		16#0a86# => X"d7e1a7e4",
		16#0a87# => X"d7e1b7e8",
		16#0a88# => X"d7e1c7ec",
		16#0a89# => X"d7e1d7f0",
		16#0a8a# => X"d7e1e7f4",
		16#0a8b# => X"d7e1f7f8",
		16#0a8c# => X"07ffff8e",
		16#0a8d# => X"9c21ff74",
		16#0a8e# => X"a860c87e",
		16#0a8f# => X"0400175c",
		16#0a90# => X"a84b0000",
		16#0a91# => X"b8820002",
		16#0a92# => X"b8420004",
		16#0a93# => X"a860c87c",
		16#0a94# => X"e2c41000",
		16#0a95# => X"18400001",
		16#0a96# => X"18800001",
		16#0a97# => X"a8426e84",
		16#0a98# => X"a8846fec",
		16#0a99# => X"e0561000",
		16#0a9a# => X"e0962000",
		16#0a9b# => X"d4025800",
		16#0a9c# => X"d4012004",
		16#0a9d# => X"0400174e",
		16#0a9e# => X"d4011000",
		16#0a9f# => X"9d6b0001",
		16#0aa0# => X"a860c87d",
		16#0aa1# => X"9ca20010",
		16#0aa2# => X"d4025804",
		16#0aa3# => X"04001748",
		16#0aa4# => X"d4012824",
		16#0aa5# => X"9d6b0001",
		16#0aa6# => X"a860c87f",
		16#0aa7# => X"d402580c",
		16#0aa8# => X"04001743",
		16#0aa9# => X"9e020008",
		16#0aaa# => X"84c10004",
		16#0aab# => X"84410024",
		16#0aac# => X"9cc60010",
		16#0aad# => X"a86b0000",
		16#0aae# => X"d4025800",
		16#0aaf# => X"04000c1c",
		16#0ab0# => X"d4013028",
		16#0ab1# => X"84810000",
		16#0ab2# => X"84a10004",
		16#0ab3# => X"84640000",
		16#0ab4# => X"9dc50008",
		16#0ab5# => X"04000c16",
		16#0ab6# => X"aa4b0000",
		16#0ab7# => X"18c00001",
		16#0ab8# => X"a88b0000",
		16#0ab9# => X"a8c670a0",
		16#0aba# => X"a8720000",
		16#0abb# => X"04000a65",
		16#0abc# => X"e3d63000",
		16#0abd# => X"a860c8be",
		16#0abe# => X"d4105800",
		16#0abf# => X"0400172c",
		16#0ac0# => X"9e5e0008",
		16#0ac1# => X"84410004",
		16#0ac2# => X"a860c8bc",
		16#0ac3# => X"04001728",
		16#0ac4# => X"d4025800",
		16#0ac5# => X"9d6b0001",
		16#0ac6# => X"a860c8bd",
		16#0ac7# => X"9c9e0010",
		16#0ac8# => X"d4025804",
		16#0ac9# => X"04001722",
		16#0aca# => X"d401202c",
		16#0acb# => X"9d6b0001",
		16#0acc# => X"a860c8bf",
		16#0acd# => X"0400171e",
		16#0ace# => X"d402580c",
		16#0acf# => X"18a00001",
		16#0ad0# => X"84c10028",
		16#0ad1# => X"a8a57154",
		16#0ad2# => X"d4065800",
		16#0ad3# => X"a86b0000",
		16#0ad4# => X"04000bf7",
		16#0ad5# => X"e3962800",
		16#0ad6# => X"84620000",
		16#0ad7# => X"9c5c0010",
		16#0ad8# => X"aa0b0000",
		16#0ad9# => X"04000bf2",
		16#0ada# => X"d4011030",
		16#0adb# => X"a8700000",
		16#0adc# => X"a88b0000",
		16#0add# => X"04000a43",
		16#0ade# => X"18400001",
		16#0adf# => X"a860c8fe",
		16#0ae0# => X"d40e5800",
		16#0ae1# => X"0400170a",
		16#0ae2# => X"a84272bc",
		16#0ae3# => X"a860c8fc",
		16#0ae4# => X"d41e5800",
		16#0ae5# => X"04001706",
		16#0ae6# => X"e3161000",
		16#0ae7# => X"18800001",
		16#0ae8# => X"9d6b0001",
		16#0ae9# => X"a860c8fd",
		16#0aea# => X"a8847208",
		16#0aeb# => X"d41e5804",
		16#0aec# => X"040016ff",
		16#0aed# => X"e3562000",
		16#0aee# => X"9d6b0001",
		16#0aef# => X"a860c8ff",
		16#0af0# => X"9cba0010",
		16#0af1# => X"d41e580c",
		16#0af2# => X"040016f9",
		16#0af3# => X"d4012834",
		16#0af4# => X"84c1002c",
		16#0af5# => X"a86b0000",
		16#0af6# => X"d4065800",
		16#0af7# => X"04000bd4",
		16#0af8# => X"9e1c0008",
		16#0af9# => X"847e0000",
		16#0afa# => X"04000bd1",
		16#0afb# => X"aa8b0000",
		16#0afc# => X"9cb80010",
		16#0afd# => X"a88b0000",
		16#0afe# => X"a8740000",
		16#0aff# => X"04000a21",
		16#0b00# => X"d4012838",
		16#0b01# => X"a860c93e",
		16#0b02# => X"d4125800",
		16#0b03# => X"040016e8",
		16#0b04# => X"9dda0008",
		16#0b05# => X"a860c93c",
		16#0b06# => X"d41c5800",
		16#0b07# => X"040016e4",
		16#0b08# => X"9c580008",
		16#0b09# => X"9d6b0001",
		16#0b0a# => X"a860c93d",
		16#0b0b# => X"040016e0",
		16#0b0c# => X"d41c5804",
		16#0b0d# => X"18c00001",
		16#0b0e# => X"9d6b0001",
		16#0b0f# => X"a8c67370",
		16#0b10# => X"a860c93f",
		16#0b11# => X"d41c580c",
		16#0b12# => X"040016d9",
		16#0b13# => X"e2963000",
		16#0b14# => X"84810030",
		16#0b15# => X"9c740010",
		16#0b16# => X"d4045800",
		16#0b17# => X"d401183c",
		16#0b18# => X"04000bb3",
		16#0b19# => X"a86b0000",
		16#0b1a# => X"9cb40008",
		16#0b1b# => X"847c0000",
		16#0b1c# => X"d4012820",
		16#0b1d# => X"04000bae",
		16#0b1e# => X"aa4b0000",
		16#0b1f# => X"18c00001",
		16#0b20# => X"a88b0000",
		16#0b21# => X"a8c67424",
		16#0b22# => X"a8720000",
		16#0b23# => X"040009fd",
		16#0b24# => X"e2563000",
		16#0b25# => X"a860c97e",
		16#0b26# => X"040016c5",
		16#0b27# => X"d4105800",
		16#0b28# => X"a860c97c",
		16#0b29# => X"040016c2",
		16#0b2a# => X"d41a5800",
		16#0b2b# => X"9d6b0001",
		16#0b2c# => X"a860c97d",
		16#0b2d# => X"9c920008",
		16#0b2e# => X"d41a5804",
		16#0b2f# => X"040016bc",
		16#0b30# => X"d4012040",
		16#0b31# => X"18a00001",
		16#0b32# => X"9d6b0001",
		16#0b33# => X"a8a57910",
		16#0b34# => X"a860c97f",
		16#0b35# => X"e0b62800",
		16#0b36# => X"d41a580c",
		16#0b37# => X"040016b4",
		16#0b38# => X"d4012808",
		16#0b39# => X"84810034",
		16#0b3a# => X"84c10008",
		16#0b3b# => X"d4045800",
		16#0b3c# => X"9cc60008",
		16#0b3d# => X"a86b0000",
		16#0b3e# => X"04000b8d",
		16#0b3f# => X"d4013044",
		16#0b40# => X"18a00001",
		16#0b41# => X"847a0000",
		16#0b42# => X"a8a579c4",
		16#0b43# => X"aa0b0000",
		16#0b44# => X"e0b62800",
		16#0b45# => X"04000b86",
		16#0b46# => X"d401280c",
		16#0b47# => X"84c1000c",
		16#0b48# => X"a88b0000",
		16#0b49# => X"9cc60008",
		16#0b4a# => X"a8700000",
		16#0b4b# => X"040009d5",
		16#0b4c# => X"d4013048",
		16#0b4d# => X"a860c9be",
		16#0b4e# => X"0400169d",
		16#0b4f# => X"d40e5800",
		16#0b50# => X"a860c9bc",
		16#0b51# => X"0400169a",
		16#0b52# => X"d4185800",
		16#0b53# => X"18800001",
		16#0b54# => X"9d6b0001",
		16#0b55# => X"a88474d8",
		16#0b56# => X"a860c9bd",
		16#0b57# => X"e0962000",
		16#0b58# => X"d4185804",
		16#0b59# => X"04001692",
		16#0b5a# => X"d4012010",
		16#0b5b# => X"84a10010",
		16#0b5c# => X"9d6b0001",
		16#0b5d# => X"a860c9bf",
		16#0b5e# => X"9ca50008",
		16#0b5f# => X"d418580c",
		16#0b60# => X"0400168b",
		16#0b61# => X"d401284c",
		16#0b62# => X"18c00001",
		16#0b63# => X"84810038",
		16#0b64# => X"a8c6758c",
		16#0b65# => X"d4045800",
		16#0b66# => X"e0d63000",
		16#0b67# => X"a86b0000",
		16#0b68# => X"04000b63",
		16#0b69# => X"d4013014",
		16#0b6a# => X"84a10014",
		16#0b6b# => X"84780000",
		16#0b6c# => X"9ca50008",
		16#0b6d# => X"a9cb0000",
		16#0b6e# => X"04000b5d",
		16#0b6f# => X"d4012850",
		16#0b70# => X"18c00001",
		16#0b71# => X"a88b0000",
		16#0b72# => X"a8c67640",
		16#0b73# => X"a86e0000",
		16#0b74# => X"e0d63000",
		16#0b75# => X"040009ab",
		16#0b76# => X"d4013018",
		16#0b77# => X"a860c9fe",
		16#0b78# => X"04001673",
		16#0b79# => X"d4025800",
		16#0b7a# => X"a860c9fc",
		16#0b7b# => X"04001670",
		16#0b7c# => X"d4145800",
		16#0b7d# => X"84410018",
		16#0b7e# => X"9d6b0001",
		16#0b7f# => X"a860c9fd",
		16#0b80# => X"9c420008",
		16#0b81# => X"d4145804",
		16#0b82# => X"04001669",
		16#0b83# => X"d4011054",
		16#0b84# => X"18800001",
		16#0b85# => X"9d6b0001",
		16#0b86# => X"a88476f4",
		16#0b87# => X"a860c9ff",
		16#0b88# => X"e0962000",
		16#0b89# => X"d414580c",
		16#0b8a# => X"04001661",
		16#0b8b# => X"d401201c",
		16#0b8c# => X"84c1003c",
		16#0b8d# => X"84a1001c",
		16#0b8e# => X"d4065800",
		16#0b8f# => X"9ca50008",
		16#0b90# => X"a86b0000",
		16#0b91# => X"18400001",
		16#0b92# => X"d4012858",
		16#0b93# => X"04000b38",
		16#0b94# => X"a84277a8",
		16#0b95# => X"84740000",
		16#0b96# => X"e2161000",
		16#0b97# => X"04000b34",
		16#0b98# => X"a9cb0000",
		16#0b99# => X"9cb00008",
		16#0b9a# => X"a88b0000",
		16#0b9b# => X"a86e0000",
		16#0b9c# => X"04000984",
		16#0b9d# => X"d401285c",
		16#0b9e# => X"84c10020",
		16#0b9f# => X"a860ca3e",
		16#0ba0# => X"0400164b",
		16#0ba1# => X"d4065800",
		16#0ba2# => X"a860ca3c",
		16#0ba3# => X"04001648",
		16#0ba4# => X"d4125800",
		16#0ba5# => X"18800001",
		16#0ba6# => X"9d6b0001",
		16#0ba7# => X"a860ca3d",
		16#0ba8# => X"a884785c",
		16#0ba9# => X"d4125804",
		16#0baa# => X"04001641",
		16#0bab# => X"e0562000",
		16#0bac# => X"9d6b0001",
		16#0bad# => X"a860ca3f",
		16#0bae# => X"9ca20008",
		16#0baf# => X"d412580c",
		16#0bb0# => X"0400163b",
		16#0bb1# => X"d4012820",
		16#0bb2# => X"a86b0000",
		16#0bb3# => X"04000b18",
		16#0bb4# => X"d4125810",
		16#0bb5# => X"84720000",
		16#0bb6# => X"04000b15",
		16#0bb7# => X"a9cb0000",
		16#0bb8# => X"a86e0000",
		16#0bb9# => X"04000967",
		16#0bba# => X"a88b0000",
		16#0bbb# => X"84c10040",
		16#0bbc# => X"a860ca7e",
		16#0bbd# => X"0400162e",
		16#0bbe# => X"d4065800",
		16#0bbf# => X"84810008",
		16#0bc0# => X"a860ca7c",
		16#0bc1# => X"0400162a",
		16#0bc2# => X"d4045800",
		16#0bc3# => X"84a10008",
		16#0bc4# => X"9d6b0001",
		16#0bc5# => X"a860ca7d",
		16#0bc6# => X"04001625",
		16#0bc7# => X"d4055804",
		16#0bc8# => X"84c10008",
		16#0bc9# => X"9d6b0001",
		16#0bca# => X"a860ca7f",
		16#0bcb# => X"04001620",
		16#0bcc# => X"d406580c",
		16#0bcd# => X"84810008",
		16#0bce# => X"a86b0000",
		16#0bcf# => X"04000afc",
		16#0bd0# => X"d4045810",
		16#0bd1# => X"84a10008",
		16#0bd2# => X"a9cb0000",
		16#0bd3# => X"04000af8",
		16#0bd4# => X"84650000",
		16#0bd5# => X"a86e0000",
		16#0bd6# => X"0400094a",
		16#0bd7# => X"a88b0000",
		16#0bd8# => X"84c10044",
		16#0bd9# => X"a860cabe",
		16#0bda# => X"04001611",
		16#0bdb# => X"d4065800",
		16#0bdc# => X"8481000c",
		16#0bdd# => X"a860cabc",
		16#0bde# => X"0400160d",
		16#0bdf# => X"d4045800",
		16#0be0# => X"84a1000c",
		16#0be1# => X"9d6b0001",
		16#0be2# => X"a860cabd",
		16#0be3# => X"04001608",
		16#0be4# => X"d4055804",
		16#0be5# => X"84c1000c",
		16#0be6# => X"9d6b0001",
		16#0be7# => X"a860cabf",
		16#0be8# => X"04001603",
		16#0be9# => X"d406580c",
		16#0bea# => X"8481000c",
		16#0beb# => X"a86b0000",
		16#0bec# => X"04000adf",
		16#0bed# => X"d4045810",
		16#0bee# => X"84a1000c",
		16#0bef# => X"a9cb0000",
		16#0bf0# => X"04000adb",
		16#0bf1# => X"84650000",
		16#0bf2# => X"a86e0000",
		16#0bf3# => X"0400092d",
		16#0bf4# => X"a88b0000",
		16#0bf5# => X"84c10048",
		16#0bf6# => X"a860cafe",
		16#0bf7# => X"040015f4",
		16#0bf8# => X"d4065800",
		16#0bf9# => X"84810010",
		16#0bfa# => X"a860cafc",
		16#0bfb# => X"040015f0",
		16#0bfc# => X"d4045800",
		16#0bfd# => X"84a10010",
		16#0bfe# => X"9d6b0001",
		16#0bff# => X"a860cafd",
		16#0c00# => X"040015eb",
		16#0c01# => X"d4055804",
		16#0c02# => X"84c10010",
		16#0c03# => X"9d6b0001",
		16#0c04# => X"a860caff",
		16#0c05# => X"040015e6",
		16#0c06# => X"d406580c",
		16#0c07# => X"84810010",
		16#0c08# => X"a86b0000",
		16#0c09# => X"04000ac2",
		16#0c0a# => X"d4045810",
		16#0c0b# => X"84a10010",
		16#0c0c# => X"a9cb0000",
		16#0c0d# => X"04000abe",
		16#0c0e# => X"84650000",
		16#0c0f# => X"a86e0000",
		16#0c10# => X"04000910",
		16#0c11# => X"a88b0000",
		16#0c12# => X"84c1004c",
		16#0c13# => X"a860cb3e",
		16#0c14# => X"040015d7",
		16#0c15# => X"d4065800",
		16#0c16# => X"84810014",
		16#0c17# => X"a860cb3c",
		16#0c18# => X"040015d3",
		16#0c19# => X"d4045800",
		16#0c1a# => X"84a10014",
		16#0c1b# => X"9d6b0001",
		16#0c1c# => X"a860cb3d",
		16#0c1d# => X"040015ce",
		16#0c1e# => X"d4055804",
		16#0c1f# => X"84c10014",
		16#0c20# => X"9d6b0001",
		16#0c21# => X"a860cb3f",
		16#0c22# => X"040015c9",
		16#0c23# => X"d406580c",
		16#0c24# => X"84810014",
		16#0c25# => X"a86b0000",
		16#0c26# => X"04000aa5",
		16#0c27# => X"d4045810",
		16#0c28# => X"84a10014",
		16#0c29# => X"a9cb0000",
		16#0c2a# => X"04000aa1",
		16#0c2b# => X"84650000",
		16#0c2c# => X"a86e0000",
		16#0c2d# => X"040008f3",
		16#0c2e# => X"a88b0000",
		16#0c2f# => X"84c10050",
		16#0c30# => X"a860cb7e",
		16#0c31# => X"040015ba",
		16#0c32# => X"d4065800",
		16#0c33# => X"84810018",
		16#0c34# => X"a860cb7c",
		16#0c35# => X"040015b6",
		16#0c36# => X"d4045800",
		16#0c37# => X"84a10018",
		16#0c38# => X"9d6b0001",
		16#0c39# => X"a860cb7d",
		16#0c3a# => X"040015b1",
		16#0c3b# => X"d4055804",
		16#0c3c# => X"84c10018",
		16#0c3d# => X"9d6b0001",
		16#0c3e# => X"a860cb7f",
		16#0c3f# => X"040015ac",
		16#0c40# => X"d406580c",
		16#0c41# => X"84810018",
		16#0c42# => X"a86b0000",
		16#0c43# => X"04000a88",
		16#0c44# => X"d4045810",
		16#0c45# => X"84a10018",
		16#0c46# => X"a9cb0000",
		16#0c47# => X"04000a84",
		16#0c48# => X"84650000",
		16#0c49# => X"a86e0000",
		16#0c4a# => X"040008d6",
		16#0c4b# => X"a88b0000",
		16#0c4c# => X"84c10054",
		16#0c4d# => X"a860cbbe",
		16#0c4e# => X"0400159d",
		16#0c4f# => X"d4065800",
		16#0c50# => X"8481001c",
		16#0c51# => X"a860cbbc",
		16#0c52# => X"04001599",
		16#0c53# => X"d4045800",
		16#0c54# => X"84a1001c",
		16#0c55# => X"9d6b0001",
		16#0c56# => X"a860cbbd",
		16#0c57# => X"04001594",
		16#0c58# => X"d4055804",
		16#0c59# => X"84c1001c",
		16#0c5a# => X"9d6b0001",
		16#0c5b# => X"a860cbbf",
		16#0c5c# => X"0400158f",
		16#0c5d# => X"d406580c",
		16#0c5e# => X"8481001c",
		16#0c5f# => X"a86b0000",
		16#0c60# => X"04000a6b",
		16#0c61# => X"d4045810",
		16#0c62# => X"84a1001c",
		16#0c63# => X"a9cb0000",
		16#0c64# => X"04000a67",
		16#0c65# => X"84650000",
		16#0c66# => X"a86e0000",
		16#0c67# => X"040008b9",
		16#0c68# => X"a88b0000",
		16#0c69# => X"84c10058",
		16#0c6a# => X"a860cbfe",
		16#0c6b# => X"04001580",
		16#0c6c# => X"d4065800",
		16#0c6d# => X"a860cbfc",
		16#0c6e# => X"0400157d",
		16#0c6f# => X"d4105800",
		16#0c70# => X"9d6b0001",
		16#0c71# => X"a860cbfd",
		16#0c72# => X"04001579",
		16#0c73# => X"d4105804",
		16#0c74# => X"9d6b0001",
		16#0c75# => X"a860cbff",
		16#0c76# => X"04001575",
		16#0c77# => X"d410580c",
		16#0c78# => X"a86b0000",
		16#0c79# => X"04000a52",
		16#0c7a# => X"d4105810",
		16#0c7b# => X"84700000",
		16#0c7c# => X"04000a4f",
		16#0c7d# => X"a9cb0000",
		16#0c7e# => X"a86e0000",
		16#0c7f# => X"040008a1",
		16#0c80# => X"a88b0000",
		16#0c81# => X"8481005c",
		16#0c82# => X"a860cc3e",
		16#0c83# => X"04001568",
		16#0c84# => X"d4045800",
		16#0c85# => X"a860cc3c",
		16#0c86# => X"04001565",
		16#0c87# => X"d4025800",
		16#0c88# => X"9d6b0001",
		16#0c89# => X"a860cc3d",
		16#0c8a# => X"04001561",
		16#0c8b# => X"d4025804",
		16#0c8c# => X"9d6b0001",
		16#0c8d# => X"a860cc3f",
		16#0c8e# => X"0400155d",
		16#0c8f# => X"d402580c",
		16#0c90# => X"a86b0000",
		16#0c91# => X"04000a3a",
		16#0c92# => X"d4025810",
		16#0c93# => X"84620000",
		16#0c94# => X"04000a37",
		16#0c95# => X"a9cb0000",
		16#0c96# => X"a86e0000",
		16#0c97# => X"04000889",
		16#0c98# => X"a88b0000",
		16#0c99# => X"84c10028",
		16#0c9a# => X"84410024",
		16#0c9b# => X"84a60000",
		16#0c9c# => X"84620000",
		16#0c9d# => X"8481002c",
		16#0c9e# => X"e0a51800",
		16#0c9f# => X"84c40000",
		16#0ca0# => X"84610004",
		16#0ca1# => X"84810000",
		16#0ca2# => X"84430000",
		16#0ca3# => X"84640000",
		16#0ca4# => X"e0a53000",
		16#0ca5# => X"e0421800",
		16#0ca6# => X"84610030",
		16#0ca7# => X"84810034",
		16#0ca8# => X"84c30000",
		16#0ca9# => X"847e0000",
		16#0caa# => X"e0a53000",
		16#0cab# => X"e0421800",
		16#0cac# => X"847c0000",
		16#0cad# => X"84c40000",
		16#0cae# => X"e0421800",
		16#0caf# => X"84610038",
		16#0cb0# => X"8481003c",
		16#0cb1# => X"e0a53000",
		16#0cb2# => X"84c30000",
		16#0cb3# => X"847a0000",
		16#0cb4# => X"e0a53000",
		16#0cb5# => X"84c40000",
		16#0cb6# => X"e0421800",
		16#0cb7# => X"e0a53000",
		16#0cb8# => X"84780000",
		16#0cb9# => X"18c00001",
		16#0cba# => X"e0421800",
		16#0cbb# => X"a8c66f38",
		16#0cbc# => X"84740000",
		16#0cbd# => X"e0963000",
		16#0cbe# => X"e0421800",
		16#0cbf# => X"84c10020",
		16#0cc0# => X"a8650000",
		16#0cc1# => X"d4042810",
		16#0cc2# => X"d4041000",
		16#0cc3# => X"d4065800",
		16#0cc4# => X"04000a07",
		16#0cc5# => X"9dc40008",
		16#0cc6# => X"a8620000",
		16#0cc7# => X"04000a04",
		16#0cc8# => X"aa0b0000",
		16#0cc9# => X"a8700000",
		16#0cca# => X"04000856",
		16#0ccb# => X"a88b0000",
		16#0ccc# => X"d40e5800",
		16#0ccd# => X"9c21008c",
		16#0cce# => X"8521fffc",
		16#0ccf# => X"8441ffd4",
		16#0cd0# => X"85c1ffd8",
		16#0cd1# => X"8601ffdc",
		16#0cd2# => X"8641ffe0",
		16#0cd3# => X"8681ffe4",
		16#0cd4# => X"86c1ffe8",
		16#0cd5# => X"8701ffec",
		16#0cd6# => X"8741fff0",
		16#0cd7# => X"8781fff4",
		16#0cd8# => X"44004800",
		16#0cd9# => X"87c1fff8",
		16#0cda# => X"d7e14ffc",
		16#0cdb# => X"d7e117d4",
		16#0cdc# => X"d7e177d8",
		16#0cdd# => X"d7e187dc",
		16#0cde# => X"d7e197e0",
		16#0cdf# => X"d7e1a7e4",
		16#0ce0# => X"d7e1b7e8",
		16#0ce1# => X"d7e1c7ec",
		16#0ce2# => X"d7e1d7f0",
		16#0ce3# => X"d7e1e7f4",
		16#0ce4# => X"d7e1f7f8",
		16#0ce5# => X"07fffd35",
		16#0ce6# => X"9c21ff98",
		16#0ce7# => X"18600001",
		16#0ce8# => X"a84b0000",
		16#0ce9# => X"a8633b09",
		16#0cea# => X"04001564",
		16#0ceb# => X"d4015800",
		16#0cec# => X"18600001",
		16#0ced# => X"d4011000",
		16#0cee# => X"a8633b55",
		16#0cef# => X"0400155f",
		16#0cf0# => X"b9c20002",
		16#0cf1# => X"18800001",
		16#0cf2# => X"18600001",
		16#0cf3# => X"a8843b9f",
		16#0cf4# => X"a8633b79",
		16#0cf5# => X"d4012004",
		16#0cf6# => X"18800001",
		16#0cf7# => X"d4011000",
		16#0cf8# => X"a8843ba5",
		16#0cf9# => X"d4012008",
		16#0cfa# => X"18800001",
		16#0cfb# => X"a8843bab",
		16#0cfc# => X"d401200c",
		16#0cfd# => X"18800001",
		16#0cfe# => X"a8843baf",
		16#0cff# => X"d4012010",
		16#0d00# => X"18800001",
		16#0d01# => X"a8843bb3",
		16#0d02# => X"d4012014",
		16#0d03# => X"18800001",
		16#0d04# => X"a8843bb7",
		16#0d05# => X"d4012018",
		16#0d06# => X"18800001",
		16#0d07# => X"a8843bbd",
		16#0d08# => X"04001546",
		16#0d09# => X"d401201c",
		16#0d0a# => X"18600001",
		16#0d0b# => X"d4011000",
		16#0d0c# => X"04001542",
		16#0d0d# => X"a8633b09",
		16#0d0e# => X"b8620004",
		16#0d0f# => X"18800001",
		16#0d10# => X"d4011000",
		16#0d11# => X"e1ce1800",
		16#0d12# => X"18600001",
		16#0d13# => X"a8846f38",
		16#0d14# => X"a8633bec",
		16#0d15# => X"e08e2000",
		16#0d16# => X"d4011804",
		16#0d17# => X"18600001",
		16#0d18# => X"d4012030",
		16#0d19# => X"a8636e84",
		16#0d1a# => X"e20e1800",
		16#0d1b# => X"84700008",
		16#0d1c# => X"84b00000",
		16#0d1d# => X"84900004",
		16#0d1e# => X"86500010",
		16#0d1f# => X"d4012808",
		16#0d20# => X"04000a38",
		16#0d21# => X"d401200c",
		16#0d22# => X"8490000c",
		16#0d23# => X"84a10030",
		16#0d24# => X"a8720000",
		16#0d25# => X"9ec50010",
		16#0d26# => X"d4015810",
		16#0d27# => X"d4016014",
		16#0d28# => X"d4012018",
		16#0d29# => X"040009a2",
		16#0d2a# => X"d401901c",
		16#0d2b# => X"18c00001",
		16#0d2c# => X"84760000",
		16#0d2d# => X"a8c66fec",
		16#0d2e# => X"aa4b0000",
		16#0d2f# => X"0400099c",
		16#0d30# => X"e20e3000",
		16#0d31# => X"18a00001",
		16#0d32# => X"a88b0000",
		16#0d33# => X"a8a570a0",
		16#0d34# => X"a8720000",
		16#0d35# => X"040007eb",
		16#0d36# => X"e28e2800",
		16#0d37# => X"18c00001",
		16#0d38# => X"a86b0000",
		16#0d39# => X"a8c67154",
		16#0d3a# => X"04000a1e",
		16#0d3b# => X"e24e3000",
		16#0d3c# => X"18600001",
		16#0d3d# => X"d4015820",
		16#0d3e# => X"d4016024",
		16#0d3f# => X"0400150f",
		16#0d40# => X"a8633bc2",
		16#0d41# => X"18800001",
		16#0d42# => X"84700008",
		16#0d43# => X"84d00000",
		16#0d44# => X"84b00004",
		16#0d45# => X"a8843bf0",
		16#0d46# => X"87100010",
		16#0d47# => X"d4013008",
		16#0d48# => X"d401280c",
		16#0d49# => X"d4011000",
		16#0d4a# => X"04000a0e",
		16#0d4b# => X"d4012004",
		16#0d4c# => X"8490000c",
		16#0d4d# => X"a8780000",
		16#0d4e# => X"d4015810",
		16#0d4f# => X"d4016014",
		16#0d50# => X"d4012018",
		16#0d51# => X"0400097a",
		16#0d52# => X"d401c01c",
		16#0d53# => X"18800001",
		16#0d54# => X"84760000",
		16#0d55# => X"a8847208",
		16#0d56# => X"ab0b0000",
		16#0d57# => X"04000974",
		16#0d58# => X"e20e2000",
		16#0d59# => X"18a00001",
		16#0d5a# => X"a88b0000",
		16#0d5b# => X"a8a572bc",
		16#0d5c# => X"a8780000",
		16#0d5d# => X"e0ae2800",
		16#0d5e# => X"040007c2",
		16#0d5f# => X"d4012828",
		16#0d60# => X"18c00001",
		16#0d61# => X"a86b0000",
		16#0d62# => X"a8c67370",
		16#0d63# => X"e0ce3000",
		16#0d64# => X"040009f4",
		16#0d65# => X"d4013034",
		16#0d66# => X"18600001",
		16#0d67# => X"d4015820",
		16#0d68# => X"d4016024",
		16#0d69# => X"040014e5",
		16#0d6a# => X"a8633bc2",
		16#0d6b# => X"18800001",
		16#0d6c# => X"84740008",
		16#0d6d# => X"84d40000",
		16#0d6e# => X"84b40004",
		16#0d6f# => X"a8843bf6",
		16#0d70# => X"87140010",
		16#0d71# => X"d4013008",
		16#0d72# => X"d401280c",
		16#0d73# => X"d4011000",
		16#0d74# => X"040009e4",
		16#0d75# => X"d4012004",
		16#0d76# => X"8494000c",
		16#0d77# => X"a8780000",
		16#0d78# => X"d4015810",
		16#0d79# => X"d4016014",
		16#0d7a# => X"d4012018",
		16#0d7b# => X"04000950",
		16#0d7c# => X"d401c01c",
		16#0d7d# => X"18800001",
		16#0d7e# => X"84760000",
		16#0d7f# => X"a8847424",
		16#0d80# => X"ab0b0000",
		16#0d81# => X"0400094a",
		16#0d82# => X"e28e2000",
		16#0d83# => X"18a00001",
		16#0d84# => X"a88b0000",
		16#0d85# => X"a8a574d8",
		16#0d86# => X"a8780000",
		16#0d87# => X"e0ae2800",
		16#0d88# => X"04000798",
		16#0d89# => X"d4012838",
		16#0d8a# => X"18c00001",
		16#0d8b# => X"a86b0000",
		16#0d8c# => X"a8c6758c",
		16#0d8d# => X"040009cb",
		16#0d8e# => X"e3ce3000",
		16#0d8f# => X"18600001",
		16#0d90# => X"d4015820",
		16#0d91# => X"d4016024",
		16#0d92# => X"040014bc",
		16#0d93# => X"a8633bc2",
		16#0d94# => X"18800001",
		16#0d95# => X"84720008",
		16#0d96# => X"84d20000",
		16#0d97# => X"84b20004",
		16#0d98# => X"a8843d68",
		16#0d99# => X"87120010",
		16#0d9a# => X"d4013008",
		16#0d9b# => X"d401280c",
		16#0d9c# => X"d4011000",
		16#0d9d# => X"040009bb",
		16#0d9e# => X"d4012004",
		16#0d9f# => X"8492000c",
		16#0da0# => X"a8780000",
		16#0da1# => X"d4015810",
		16#0da2# => X"d4016014",
		16#0da3# => X"d4012018",
		16#0da4# => X"04000927",
		16#0da5# => X"d401c01c",
		16#0da6# => X"18800001",
		16#0da7# => X"84760000",
		16#0da8# => X"a8847640",
		16#0da9# => X"ab0b0000",
		16#0daa# => X"04000921",
		16#0dab# => X"e38e2000",
		16#0dac# => X"18a00001",
		16#0dad# => X"a88b0000",
		16#0dae# => X"a8a576f4",
		16#0daf# => X"a8780000",
		16#0db0# => X"04000770",
		16#0db1# => X"e34e2800",
		16#0db2# => X"18c00001",
		16#0db3# => X"a86b0000",
		16#0db4# => X"a8c677a8",
		16#0db5# => X"040009a3",
		16#0db6# => X"e30e3000",
		16#0db7# => X"18600001",
		16#0db8# => X"d4015820",
		16#0db9# => X"d4016024",
		16#0dba# => X"04001494",
		16#0dbb# => X"a8633bc2",
		16#0dbc# => X"18800001",
		16#0dbd# => X"84700008",
		16#0dbe# => X"84d00000",
		16#0dbf# => X"84b00004",
		16#0dc0# => X"a8843d72",
		16#0dc1# => X"d4013008",
		16#0dc2# => X"d401280c",
		16#0dc3# => X"d4011000",
		16#0dc4# => X"04000994",
		16#0dc5# => X"d4012004",
		16#0dc6# => X"8490000c",
		16#0dc7# => X"84700010",
		16#0dc8# => X"d4015810",
		16#0dc9# => X"d4016014",
		16#0dca# => X"d4012018",
		16#0dcb# => X"04000900",
		16#0dcc# => X"d401181c",
		16#0dcd# => X"18a00001",
		16#0dce# => X"84760000",
		16#0dcf# => X"a8a5785c",
		16#0dd0# => X"d401582c",
		16#0dd1# => X"040008fa",
		16#0dd2# => X"e1ce2800",
		16#0dd3# => X"8461002c",
		16#0dd4# => X"0400074c",
		16#0dd5# => X"a88b0000",
		16#0dd6# => X"04000982",
		16#0dd7# => X"a86b0000",
		16#0dd8# => X"18600001",
		16#0dd9# => X"d4015820",
		16#0dda# => X"d4016024",
		16#0ddb# => X"04001473",
		16#0ddc# => X"a8633bc2",
		16#0ddd# => X"84810028",
		16#0dde# => X"84c10028",
		16#0ddf# => X"84a40004",
		16#0de0# => X"84840010",
		16#0de1# => X"84660008",
		16#0de2# => X"84c60000",
		16#0de3# => X"d401201c",
		16#0de4# => X"18800001",
		16#0de5# => X"d4013008",
		16#0de6# => X"a8843bfa",
		16#0de7# => X"d4011000",
		16#0de8# => X"d4012004",
		16#0de9# => X"0400096f",
		16#0dea# => X"d401280c",
		16#0deb# => X"84a10028",
		16#0dec# => X"8461001c",
		16#0ded# => X"8485000c",
		16#0dee# => X"d4015810",
		16#0def# => X"d4016014",
		16#0df0# => X"040008db",
		16#0df1# => X"d4012018",
		16#0df2# => X"84760000",
		16#0df3# => X"040008d8",
		16#0df4# => X"d4015828",
		16#0df5# => X"84610028",
		16#0df6# => X"0400072a",
		16#0df7# => X"a88b0000",
		16#0df8# => X"04000960",
		16#0df9# => X"a86b0000",
		16#0dfa# => X"18600001",
		16#0dfb# => X"d4015820",
		16#0dfc# => X"d4016024",
		16#0dfd# => X"04001451",
		16#0dfe# => X"a8633bc2",
		16#0dff# => X"84810034",
		16#0e00# => X"84c10034",
		16#0e01# => X"84a40004",
		16#0e02# => X"84840010",
		16#0e03# => X"84660008",
		16#0e04# => X"84c60000",
		16#0e05# => X"d401201c",
		16#0e06# => X"18800001",
		16#0e07# => X"d4013008",
		16#0e08# => X"a8843bff",
		16#0e09# => X"d4011000",
		16#0e0a# => X"d4012004",
		16#0e0b# => X"0400094d",
		16#0e0c# => X"d401280c",
		16#0e0d# => X"84a10034",
		16#0e0e# => X"8461001c",
		16#0e0f# => X"8485000c",
		16#0e10# => X"d4015810",
		16#0e11# => X"d4016014",
		16#0e12# => X"040008b9",
		16#0e13# => X"d4012018",
		16#0e14# => X"84760000",
		16#0e15# => X"040008b6",
		16#0e16# => X"d4015828",
		16#0e17# => X"84610028",
		16#0e18# => X"04000708",
		16#0e19# => X"a88b0000",
		16#0e1a# => X"0400093e",
		16#0e1b# => X"a86b0000",
		16#0e1c# => X"18600001",
		16#0e1d# => X"d4015820",
		16#0e1e# => X"d4016024",
		16#0e1f# => X"0400142f",
		16#0e20# => X"a8633bc2",
		16#0e21# => X"84810030",
		16#0e22# => X"84c10030",
		16#0e23# => X"84a40004",
		16#0e24# => X"18800001",
		16#0e25# => X"84660008",
		16#0e26# => X"a8843c29",
		16#0e27# => X"84c60000",
		16#0e28# => X"d4011000",
		16#0e29# => X"d4012004",
		16#0e2a# => X"d4013008",
		16#0e2b# => X"0400092d",
		16#0e2c# => X"d401280c",
		16#0e2d# => X"84c10030",
		16#0e2e# => X"18600001",
		16#0e2f# => X"84a6000c",
		16#0e30# => X"84960000",
		16#0e31# => X"a8633c05",
		16#0e32# => X"d4015810",
		16#0e33# => X"d4016014",
		16#0e34# => X"d4012818",
		16#0e35# => X"04001419",
		16#0e36# => X"d401201c",
		16#0e37# => X"18800001",
		16#0e38# => X"84740008",
		16#0e39# => X"84d40000",
		16#0e3a# => X"84b40004",
		16#0e3b# => X"a8843c30",
		16#0e3c# => X"d4013008",
		16#0e3d# => X"d4011000",
		16#0e3e# => X"d4012004",
		16#0e3f# => X"04000919",
		16#0e40# => X"d401280c",
		16#0e41# => X"18600001",
		16#0e42# => X"84b4000c",
		16#0e43# => X"84940010",
		16#0e44# => X"a8633c05",
		16#0e45# => X"d4015810",
		16#0e46# => X"d4016014",
		16#0e47# => X"d4012818",
		16#0e48# => X"04001406",
		16#0e49# => X"d401201c",
		16#0e4a# => X"84810038",
		16#0e4b# => X"84640008",
		16#0e4c# => X"86c40000",
		16#0e4d# => X"84a40004",
		16#0e4e# => X"18800001",
		16#0e4f# => X"d4011000",
		16#0e50# => X"a8843c2d",
		16#0e51# => X"d401b008",
		16#0e52# => X"d4012004",
		16#0e53# => X"04000905",
		16#0e54# => X"d401280c",
		16#0e55# => X"84c10038",
		16#0e56# => X"a8760000",
		16#0e57# => X"84a6000c",
		16#0e58# => X"84860010",
		16#0e59# => X"d4012818",
		16#0e5a# => X"d4015810",
		16#0e5b# => X"d4016014",
		16#0e5c# => X"0400086f",
		16#0e5d# => X"d401201c",
		16#0e5e# => X"84740000",
		16#0e5f# => X"0400086c",
		16#0e60# => X"aacb0000",
		16#0e61# => X"a8760000",
		16#0e62# => X"040006be",
		16#0e63# => X"a88b0000",
		16#0e64# => X"040008f4",
		16#0e65# => X"a86b0000",
		16#0e66# => X"18600001",
		16#0e67# => X"d4015820",
		16#0e68# => X"d4016024",
		16#0e69# => X"040013e5",
		16#0e6a# => X"a8633bc2",
		16#0e6b# => X"18800001",
		16#0e6c# => X"847e0008",
		16#0e6d# => X"86de0000",
		16#0e6e# => X"84be0004",
		16#0e6f# => X"a8843c34",
		16#0e70# => X"d4011000",
		16#0e71# => X"d4012004",
		16#0e72# => X"d401b008",
		16#0e73# => X"040008e5",
		16#0e74# => X"d401280c",
		16#0e75# => X"84be000c",
		16#0e76# => X"849e0010",
		16#0e77# => X"a8760000",
		16#0e78# => X"d4012818",
		16#0e79# => X"d4015810",
		16#0e7a# => X"d4016014",
		16#0e7b# => X"04000850",
		16#0e7c# => X"d401201c",
		16#0e7d# => X"84740000",
		16#0e7e# => X"0400084d",
		16#0e7f# => X"aacb0000",
		16#0e80# => X"a8760000",
		16#0e81# => X"0400069f",
		16#0e82# => X"a88b0000",
		16#0e83# => X"040008d5",
		16#0e84# => X"a86b0000",
		16#0e85# => X"18600001",
		16#0e86# => X"d4015820",
		16#0e87# => X"d4016024",
		16#0e88# => X"040013c6",
		16#0e89# => X"a8633bc2",
		16#0e8a# => X"18800001",
		16#0e8b# => X"847c0008",
		16#0e8c# => X"869c0000",
		16#0e8d# => X"84bc0004",
		16#0e8e# => X"a8843c3b",
		16#0e8f# => X"d4011000",
		16#0e90# => X"d4012004",
		16#0e91# => X"d401a008",
		16#0e92# => X"040008c6",
		16#0e93# => X"d401280c",
		16#0e94# => X"84bc000c",
		16#0e95# => X"849c0010",
		16#0e96# => X"a8740000",
		16#0e97# => X"d4012818",
		16#0e98# => X"d4015810",
		16#0e99# => X"d4016014",
		16#0e9a# => X"04000831",
		16#0e9b# => X"d401201c",
		16#0e9c# => X"84720000",
		16#0e9d# => X"0400082e",
		16#0e9e# => X"aa8b0000",
		16#0e9f# => X"a8740000",
		16#0ea0# => X"04000680",
		16#0ea1# => X"a88b0000",
		16#0ea2# => X"040008b6",
		16#0ea3# => X"a86b0000",
		16#0ea4# => X"18600001",
		16#0ea5# => X"d4015820",
		16#0ea6# => X"d4016024",
		16#0ea7# => X"040013a7",
		16#0ea8# => X"a8633bc2",
		16#0ea9# => X"18800001",
		16#0eaa# => X"847a0008",
		16#0eab# => X"869a0000",
		16#0eac# => X"84ba0004",
		16#0ead# => X"a8843c42",
		16#0eae# => X"d4011000",
		16#0eaf# => X"d4012004",
		16#0eb0# => X"d401a008",
		16#0eb1# => X"040008a7",
		16#0eb2# => X"d401280c",
		16#0eb3# => X"84ba000c",
		16#0eb4# => X"849a0010",
		16#0eb5# => X"a8740000",
		16#0eb6# => X"d4012818",
		16#0eb7# => X"d4015810",
		16#0eb8# => X"d4016014",
		16#0eb9# => X"04000812",
		16#0eba# => X"d401201c",
		16#0ebb# => X"84720000",
		16#0ebc# => X"0400080f",
		16#0ebd# => X"aa8b0000",
		16#0ebe# => X"a8740000",
		16#0ebf# => X"04000661",
		16#0ec0# => X"a88b0000",
		16#0ec1# => X"04000897",
		16#0ec2# => X"a86b0000",
		16#0ec3# => X"18600001",
		16#0ec4# => X"d4015820",
		16#0ec5# => X"d4016024",
		16#0ec6# => X"04001388",
		16#0ec7# => X"a8633bc2",
		16#0ec8# => X"18800001",
		16#0ec9# => X"84780008",
		16#0eca# => X"86580000",
		16#0ecb# => X"84b80004",
		16#0ecc# => X"a8843c49",
		16#0ecd# => X"d4011000",
		16#0ece# => X"d4012004",
		16#0ecf# => X"d4019008",
		16#0ed0# => X"04000888",
		16#0ed1# => X"d401280c",
		16#0ed2# => X"84b8000c",
		16#0ed3# => X"84980010",
		16#0ed4# => X"a8720000",
		16#0ed5# => X"d4012818",
		16#0ed6# => X"d4015810",
		16#0ed7# => X"d4016014",
		16#0ed8# => X"040007f3",
		16#0ed9# => X"d401201c",
		16#0eda# => X"84700000",
		16#0edb# => X"040007f0",
		16#0edc# => X"aa4b0000",
		16#0edd# => X"a8720000",
		16#0ede# => X"04000642",
		16#0edf# => X"a88b0000",
		16#0ee0# => X"04000878",
		16#0ee1# => X"a86b0000",
		16#0ee2# => X"18600001",
		16#0ee3# => X"d4015820",
		16#0ee4# => X"d4016024",
		16#0ee5# => X"04001369",
		16#0ee6# => X"a8633bc2",
		16#0ee7# => X"846e0008",
		16#0ee8# => X"864e0000",
		16#0ee9# => X"848e0004",
		16#0eea# => X"d4011000",
		16#0eeb# => X"18400001",
		16#0eec# => X"d4019008",
		16#0eed# => X"a8423c50",
		16#0eee# => X"d401200c",
		16#0eef# => X"04000869",
		16#0ef0# => X"d4011004",
		16#0ef1# => X"848e000c",
		16#0ef2# => X"844e0010",
		16#0ef3# => X"a8720000",
		16#0ef4# => X"d4015810",
		16#0ef5# => X"d4016014",
		16#0ef6# => X"d4012018",
		16#0ef7# => X"040007d4",
		16#0ef8# => X"d401101c",
		16#0ef9# => X"84700000",
		16#0efa# => X"040007d1",
		16#0efb# => X"a84b0000",
		16#0efc# => X"a8620000",
		16#0efd# => X"04000623",
		16#0efe# => X"a88b0000",
		16#0eff# => X"04000859",
		16#0f00# => X"a86b0000",
		16#0f01# => X"18600001",
		16#0f02# => X"d4015820",
		16#0f03# => X"d4016024",
		16#0f04# => X"0400134a",
		16#0f05# => X"a8633bc2",
		16#0f06# => X"9c210068",
		16#0f07# => X"8521fffc",
		16#0f08# => X"8441ffd4",
		16#0f09# => X"85c1ffd8",
		16#0f0a# => X"8601ffdc",
		16#0f0b# => X"8641ffe0",
		16#0f0c# => X"8681ffe4",
		16#0f0d# => X"86c1ffe8",
		16#0f0e# => X"8701ffec",
		16#0f0f# => X"8741fff0",
		16#0f10# => X"8781fff4",
		16#0f11# => X"44004800",
		16#0f12# => X"87c1fff8",
		16#0f13# => X"d7e177f8",
		16#0f14# => X"d7e14ffc",
		16#0f15# => X"d7e117f4",
		16#0f16# => X"9c21fff4",
		16#0f17# => X"07fffafd",
		16#0f18# => X"a9c30000",
		16#0f19# => X"bc0b0000",
		16#0f1a# => X"10000031",
		16#0f1b# => X"9ca00000",
		16#0f1c# => X"18c00fff",
		16#0f1d# => X"9c8e0004",
		16#0f1e# => X"a8c6ffff",
		16#0f1f# => X"a8450000",
		16#0f20# => X"84e40000",
		16#0f21# => X"e4a63800",
		16#0f22# => X"10000003",
		16#0f23# => X"9c420001",
		16#0f24# => X"a8c70000",
		16#0f25# => X"84e40008",
		16#0f26# => X"e4653800",
		16#0f27# => X"10000003",
		16#0f28# => X"9c840014",
		16#0f29# => X"a8a70000",
		16#0f2a# => X"e4825800",
		16#0f2b# => X"13fffff5",
		16#0f2c# => X"a86e0000",
		16#0f2d# => X"9c4e00a0",
		16#0f2e# => X"d4023004",
		16#0f2f# => X"d402280c",
		16#0f30# => X"84c20010",
		16#0f31# => X"84a20000",
		16#0f32# => X"9c800000",
		16#0f33# => X"85030010",
		16#0f34# => X"84e30000",
		16#0f35# => X"e0c64000",
		16#0f36# => X"e0a53800",
		16#0f37# => X"9c840001",
		16#0f38# => X"d4023010",
		16#0f39# => X"d4022800",
		16#0f3a# => X"e44b2000",
		16#0f3b# => X"13fffff8",
		16#0f3c# => X"9c630014",
		16#0f3d# => X"0400078e",
		16#0f3e# => X"84620010",
		16#0f3f# => X"84620000",
		16#0f40# => X"0400078b",
		16#0f41# => X"a9cb0000",
		16#0f42# => X"a86e0000",
		16#0f43# => X"040005dd",
		16#0f44# => X"a88b0000",
		16#0f45# => X"d4025808",
		16#0f46# => X"9c21000c",
		16#0f47# => X"8521fffc",
		16#0f48# => X"8441fff4",
		16#0f49# => X"44004800",
		16#0f4a# => X"85c1fff8",
		16#0f4b# => X"18600fff",
		16#0f4c# => X"9c4e00a0",
		16#0f4d# => X"a863ffff",
		16#0f4e# => X"d402580c",
		16#0f4f# => X"03ffffee",
		16#0f50# => X"d4021804",
		16#0f51# => X"18600001",
		16#0f52# => X"d7e14ffc",
		16#0f53# => X"d7e117f0",
		16#0f54# => X"d7e177f4",
		16#0f55# => X"d7e187f8",
		16#0f56# => X"a8636e84",
		16#0f57# => X"9c21fff0",
		16#0f58# => X"07ffffbb",
		16#0f59# => X"18400001",
		16#0f5a# => X"18600001",
		16#0f5b# => X"a8426f38",
		16#0f5c# => X"07ffffb7",
		16#0f5d# => X"a8636fec",
		16#0f5e# => X"18600001",
		16#0f5f# => X"07ffffb4",
		16#0f60# => X"a86370a0",
		16#0f61# => X"18600001",
		16#0f62# => X"07ffffb1",
		16#0f63# => X"a8637154",
		16#0f64# => X"18600001",
		16#0f65# => X"07ffffae",
		16#0f66# => X"a8637208",
		16#0f67# => X"18600001",
		16#0f68# => X"07ffffab",
		16#0f69# => X"a86372bc",
		16#0f6a# => X"18600001",
		16#0f6b# => X"07ffffa8",
		16#0f6c# => X"a8637370",
		16#0f6d# => X"18600001",
		16#0f6e# => X"07ffffa5",
		16#0f6f# => X"a8637424",
		16#0f70# => X"18600001",
		16#0f71# => X"07ffffa2",
		16#0f72# => X"a8637910",
		16#0f73# => X"18600001",
		16#0f74# => X"07ffff9f",
		16#0f75# => X"a86379c4",
		16#0f76# => X"18600001",
		16#0f77# => X"07ffff9c",
		16#0f78# => X"a86374d8",
		16#0f79# => X"18600001",
		16#0f7a# => X"07ffff99",
		16#0f7b# => X"a863758c",
		16#0f7c# => X"18600001",
		16#0f7d# => X"07ffff96",
		16#0f7e# => X"a8637640",
		16#0f7f# => X"18600001",
		16#0f80# => X"07ffff93",
		16#0f81# => X"a86376f4",
		16#0f82# => X"18600001",
		16#0f83# => X"07ffff90",
		16#0f84# => X"a86377a8",
		16#0f85# => X"18600001",
		16#0f86# => X"07ffff8d",
		16#0f87# => X"a863785c",
		16#0f88# => X"18c00001",
		16#0f89# => X"18800001",
		16#0f8a# => X"a8c66fec",
		16#0f8b# => X"a8846e84",
		16#0f8c# => X"18a00001",
		16#0f8d# => X"846400b0",
		16#0f8e# => X"84e600b0",
		16#0f8f# => X"a8a570a0",
		16#0f90# => X"e0e71800",
		16#0f91# => X"850500b0",
		16#0f92# => X"85c600a0",
		16#0f93# => X"18600001",
		16#0f94# => X"84c400a0",
		16#0f95# => X"84a500a0",
		16#0f96# => X"e0874000",
		16#0f97# => X"a8637154",
		16#0f98# => X"e1ce3000",
		16#0f99# => X"18e00001",
		16#0f9a# => X"850300b0",
		16#0f9b# => X"a8e77208",
		16#0f9c# => X"846300a0",
		16#0f9d# => X"e1ce2800",
		16#0f9e# => X"18c00001",
		16#0f9f# => X"e0844000",
		16#0fa0# => X"a8c672bc",
		16#0fa1# => X"850700b0",
		16#0fa2# => X"e1ce1800",
		16#0fa3# => X"18a00001",
		16#0fa4# => X"846700a0",
		16#0fa5# => X"e0844000",
		16#0fa6# => X"a8a57370",
		16#0fa7# => X"850600b0",
		16#0fa8# => X"e1ce1800",
		16#0fa9# => X"846600a0",
		16#0faa# => X"84e500b0",
		16#0fab# => X"e0844000",
		16#0fac# => X"84a500a0",
		16#0fad# => X"e1ce1800",
		16#0fae# => X"e0843800",
		16#0faf# => X"e1ce2800",
		16#0fb0# => X"a8640000",
		16#0fb1# => X"d40220b0",
		16#0fb2# => X"04000719",
		16#0fb3# => X"d40270a0",
		16#0fb4# => X"a86e0000",
		16#0fb5# => X"04000716",
		16#0fb6# => X"aa0b0000",
		16#0fb7# => X"a8700000",
		16#0fb8# => X"04000568",
		16#0fb9# => X"a88b0000",
		16#0fba# => X"d40258a8",
		16#0fbb# => X"9c210010",
		16#0fbc# => X"8521fffc",
		16#0fbd# => X"8441fff0",
		16#0fbe# => X"85c1fff4",
		16#0fbf# => X"44004800",
		16#0fc0# => X"8601fff8",
		16#0fc1# => X"18600001",
		16#0fc2# => X"d7e14ffc",
		16#0fc3# => X"d7e117d4",
		16#0fc4# => X"d7e177d8",
		16#0fc5# => X"d7e187dc",
		16#0fc6# => X"d7e197e0",
		16#0fc7# => X"d7e1a7e4",
		16#0fc8# => X"d7e1b7e8",
		16#0fc9# => X"d7e1c7ec",
		16#0fca# => X"d7e1d7f0",
		16#0fcb# => X"d7e1e7f4",
		16#0fcc# => X"d7e1f7f8",
		16#0fcd# => X"a8633c57",
		16#0fce# => X"9c21ffac",
		16#0fcf# => X"040012c2",
		16#0fd0# => X"19c00001",
		16#0fd1# => X"18600001",
		16#0fd2# => X"a9ce6e84",
		16#0fd3# => X"a8633ca1",
		16#0fd4# => X"040012bd",
		16#0fd5# => X"18400001",
		16#0fd6# => X"18800001",
		16#0fd7# => X"18600001",
		16#0fd8# => X"a8843b9f",
		16#0fd9# => X"a8633cca",
		16#0fda# => X"d4012000",
		16#0fdb# => X"18800001",
		16#0fdc# => X"a8426f38",
		16#0fdd# => X"a8843ba5",
		16#0fde# => X"1a400001",
		16#0fdf# => X"d4012004",
		16#0fe0# => X"18800001",
		16#0fe1# => X"aa526fec",
		16#0fe2# => X"a8843bab",
		16#0fe3# => X"1a800001",
		16#0fe4# => X"d4012008",
		16#0fe5# => X"18800001",
		16#0fe6# => X"aa9470a0",
		16#0fe7# => X"a8843baf",
		16#0fe8# => X"1bc00001",
		16#0fe9# => X"d401200c",
		16#0fea# => X"18800001",
		16#0feb# => X"abde7640",
		16#0fec# => X"a8843bb3",
		16#0fed# => X"1b800001",
		16#0fee# => X"d4012010",
		16#0fef# => X"18800001",
		16#0ff0# => X"ab9c76f4",
		16#0ff1# => X"a8843bb7",
		16#0ff2# => X"1b400001",
		16#0ff3# => X"d4012014",
		16#0ff4# => X"18800001",
		16#0ff5# => X"ab5a77a8",
		16#0ff6# => X"a8843bbd",
		16#0ff7# => X"1b000001",
		16#0ff8# => X"04001256",
		16#0ff9# => X"d4012018",
		16#0ffa# => X"18600001",
		16#0ffb# => X"ab18785c",
		16#0ffc# => X"04001295",
		16#0ffd# => X"a8633c57",
		16#0ffe# => X"18800001",
		16#0fff# => X"846e00a8",
		16#1000# => X"84ce00a0",
		16#1001# => X"84ae00a4",
		16#1002# => X"a8843bec",
		16#1003# => X"860e00b0",
		16#1004# => X"d4013004",
		16#1005# => X"d4012808",
		16#1006# => X"04000752",
		16#1007# => X"d4012000",
		16#1008# => X"848e00ac",
		16#1009# => X"a8700000",
		16#100a# => X"d401580c",
		16#100b# => X"d4016010",
		16#100c# => X"d4012014",
		16#100d# => X"040006be",
		16#100e# => X"d4018018",
		16#100f# => X"846200b0",
		16#1010# => X"040006bb",
		16#1011# => X"a9cb0000",
		16#1012# => X"a86e0000",
		16#1013# => X"a88b0000",
		16#1014# => X"0400050c",
		16#1015# => X"1a000001",
		16#1016# => X"a86b0000",
		16#1017# => X"04000741",
		16#1018# => X"aa107154",
		16#1019# => X"18600001",
		16#101a# => X"d401581c",
		16#101b# => X"d4016020",
		16#101c# => X"a8633cef",
		16#101d# => X"04001231",
		16#101e# => X"19c00001",
		16#101f# => X"18800001",
		16#1020# => X"847200a8",
		16#1021# => X"84d200a0",
		16#1022# => X"84b200a4",
		16#1023# => X"a8843bf0",
		16#1024# => X"86d200b0",
		16#1025# => X"d4013004",
		16#1026# => X"d4012808",
		16#1027# => X"04000731",
		16#1028# => X"d4012000",
		16#1029# => X"849200ac",
		16#102a# => X"a8760000",
		16#102b# => X"d401580c",
		16#102c# => X"d4016010",
		16#102d# => X"d4012014",
		16#102e# => X"0400069d",
		16#102f# => X"d401b018",
		16#1030# => X"846200b0",
		16#1031# => X"0400069a",
		16#1032# => X"aa4b0000",
		16#1033# => X"a8720000",
		16#1034# => X"a88b0000",
		16#1035# => X"040004eb",
		16#1036# => X"a9ce7208",
		16#1037# => X"a86b0000",
		16#1038# => X"04000720",
		16#1039# => X"1a400001",
		16#103a# => X"18600001",
		16#103b# => X"d401581c",
		16#103c# => X"d4016020",
		16#103d# => X"a8633cef",
		16#103e# => X"04001210",
		16#103f# => X"aa527424",
		16#1040# => X"18800001",
		16#1041# => X"847400a8",
		16#1042# => X"84d400a0",
		16#1043# => X"84b400a4",
		16#1044# => X"a8843bf6",
		16#1045# => X"86d400b0",
		16#1046# => X"d4013004",
		16#1047# => X"d4012808",
		16#1048# => X"04000710",
		16#1049# => X"d4012000",
		16#104a# => X"849400ac",
		16#104b# => X"a8760000",
		16#104c# => X"d401580c",
		16#104d# => X"d4016010",
		16#104e# => X"d4012014",
		16#104f# => X"0400067c",
		16#1050# => X"d401b018",
		16#1051# => X"846200b0",
		16#1052# => X"04000679",
		16#1053# => X"aa8b0000",
		16#1054# => X"a8740000",
		16#1055# => X"a88b0000",
		16#1056# => X"040004ca",
		16#1057# => X"1ac00001",
		16#1058# => X"a86b0000",
		16#1059# => X"040006ff",
		16#105a# => X"aad67910",
		16#105b# => X"18600001",
		16#105c# => X"d401581c",
		16#105d# => X"d4016020",
		16#105e# => X"040011f0",
		16#105f# => X"a8633cef",
		16#1060# => X"18800001",
		16#1061# => X"847000a8",
		16#1062# => X"84d000a0",
		16#1063# => X"84b000a4",
		16#1064# => X"a8843d68",
		16#1065# => X"869000b0",
		16#1066# => X"d4013004",
		16#1067# => X"d4012808",
		16#1068# => X"040006f0",
		16#1069# => X"d4012000",
		16#106a# => X"849000ac",
		16#106b# => X"a8740000",
		16#106c# => X"d401580c",
		16#106d# => X"d4016010",
		16#106e# => X"d4012014",
		16#106f# => X"0400065c",
		16#1070# => X"d401a018",
		16#1071# => X"846200b0",
		16#1072# => X"04000659",
		16#1073# => X"aa8b0000",
		16#1074# => X"a8740000",
		16#1075# => X"040004ab",
		16#1076# => X"a88b0000",
		16#1077# => X"040006e1",
		16#1078# => X"a86b0000",
		16#1079# => X"18600001",
		16#107a# => X"d401581c",
		16#107b# => X"d4016020",
		16#107c# => X"040011d2",
		16#107d# => X"a8633cef",
		16#107e# => X"18800001",
		16#107f# => X"846e00a8",
		16#1080# => X"84ce00a0",
		16#1081# => X"84ae00a4",
		16#1082# => X"a8843d72",
		16#1083# => X"868e00b0",
		16#1084# => X"d4013004",
		16#1085# => X"d4012808",
		16#1086# => X"040006d2",
		16#1087# => X"d4012000",
		16#1088# => X"848e00ac",
		16#1089# => X"a8740000",
		16#108a# => X"d401580c",
		16#108b# => X"d4016010",
		16#108c# => X"d4012014",
		16#108d# => X"0400063e",
		16#108e# => X"d401a018",
		16#108f# => X"846200b0",
		16#1090# => X"0400063b",
		16#1091# => X"aa8b0000",
		16#1092# => X"a8740000",
		16#1093# => X"a88b0000",
		16#1094# => X"0400048c",
		16#1095# => X"1a800001",
		16#1096# => X"a86b0000",
		16#1097# => X"040006c1",
		16#1098# => X"aa9479c4",
		16#1099# => X"18600001",
		16#109a# => X"d401581c",
		16#109b# => X"d4016020",
		16#109c# => X"040011b2",
		16#109d# => X"a8633cef",
		16#109e# => X"18800001",
		16#109f# => X"a88472bc",
		16#10a0# => X"84c400a0",
		16#10a1# => X"846400a8",
		16#10a2# => X"84a400a4",
		16#10a3# => X"848400b0",
		16#10a4# => X"d4013004",
		16#10a5# => X"d4012018",
		16#10a6# => X"18800001",
		16#10a7# => X"d4012808",
		16#10a8# => X"a8843bfa",
		16#10a9# => X"040006af",
		16#10aa# => X"d4012000",
		16#10ab# => X"18a00001",
		16#10ac# => X"84610018",
		16#10ad# => X"a8a572bc",
		16#10ae# => X"848500ac",
		16#10af# => X"d401580c",
		16#10b0# => X"d4016010",
		16#10b1# => X"0400061a",
		16#10b2# => X"d4012014",
		16#10b3# => X"846200b0",
		16#10b4# => X"04000617",
		16#10b5# => X"d4015824",
		16#10b6# => X"84610024",
		16#10b7# => X"04000469",
		16#10b8# => X"a88b0000",
		16#10b9# => X"0400069f",
		16#10ba# => X"a86b0000",
		16#10bb# => X"18600001",
		16#10bc# => X"d401581c",
		16#10bd# => X"d4016020",
		16#10be# => X"04001190",
		16#10bf# => X"a8633cef",
		16#10c0# => X"18800001",
		16#10c1# => X"a8847370",
		16#10c2# => X"84c400a0",
		16#10c3# => X"846400a8",
		16#10c4# => X"84a400a4",
		16#10c5# => X"848400b0",
		16#10c6# => X"d4013004",
		16#10c7# => X"d4012018",
		16#10c8# => X"18800001",
		16#10c9# => X"d4012808",
		16#10ca# => X"a8843bff",
		16#10cb# => X"0400068d",
		16#10cc# => X"d4012000",
		16#10cd# => X"18a00001",
		16#10ce# => X"84610018",
		16#10cf# => X"a8a57370",
		16#10d0# => X"848500ac",
		16#10d1# => X"d401580c",
		16#10d2# => X"d4016010",
		16#10d3# => X"040005f8",
		16#10d4# => X"d4012014",
		16#10d5# => X"846200b0",
		16#10d6# => X"040005f5",
		16#10d7# => X"d4015824",
		16#10d8# => X"84610024",
		16#10d9# => X"04000447",
		16#10da# => X"a88b0000",
		16#10db# => X"0400067d",
		16#10dc# => X"a86b0000",
		16#10dd# => X"18600001",
		16#10de# => X"d401581c",
		16#10df# => X"d4016020",
		16#10e0# => X"0400116e",
		16#10e1# => X"a8633cef",
		16#10e2# => X"848200a0",
		16#10e3# => X"84a200a4",
		16#10e4# => X"846200a8",
		16#10e5# => X"d4012004",
		16#10e6# => X"18800001",
		16#10e7# => X"d4012808",
		16#10e8# => X"a8843c29",
		16#10e9# => X"0400066f",
		16#10ea# => X"d4012000",
		16#10eb# => X"18600001",
		16#10ec# => X"848200ac",
		16#10ed# => X"a8633d18",
		16#10ee# => X"844200b0",
		16#10ef# => X"d401580c",
		16#10f0# => X"d4016010",
		16#10f1# => X"d4012014",
		16#10f2# => X"0400115c",
		16#10f3# => X"d4011018",
		16#10f4# => X"845200a0",
		16#10f5# => X"847200a8",
		16#10f6# => X"849200a4",
		16#10f7# => X"d4011004",
		16#10f8# => X"18400001",
		16#10f9# => X"d4012008",
		16#10fa# => X"a8423c30",
		16#10fb# => X"0400065d",
		16#10fc# => X"d4011000",
		16#10fd# => X"18600001",
		16#10fe# => X"849200ac",
		16#10ff# => X"845200b0",
		16#1100# => X"a8633d18",
		16#1101# => X"d401580c",
		16#1102# => X"d4016010",
		16#1103# => X"d4012014",
		16#1104# => X"0400114a",
		16#1105# => X"d4011018",
		16#1106# => X"18800001",
		16#1107# => X"18400001",
		16#1108# => X"a88474d8",
		16#1109# => X"a84274d8",
		16#110a# => X"84a400a4",
		16#110b# => X"18800001",
		16#110c# => X"846200a8",
		16#110d# => X"a8843c2d",
		16#110e# => X"844200a0",
		16#110f# => X"d4012000",
		16#1110# => X"d4011004",
		16#1111# => X"04000647",
		16#1112# => X"d4012808",
		16#1113# => X"18a00001",
		16#1114# => X"a8620000",
		16#1115# => X"a8a574d8",
		16#1116# => X"848500ac",
		16#1117# => X"844500b0",
		16#1118# => X"d401580c",
		16#1119# => X"d4016010",
		16#111a# => X"d4012014",
		16#111b# => X"040005b0",
		16#111c# => X"d4011018",
		16#111d# => X"847200a0",
		16#111e# => X"040005ad",
		16#111f# => X"a84b0000",
		16#1120# => X"a8620000",
		16#1121# => X"a88b0000",
		16#1122# => X"040003fe",
		16#1123# => X"18400001",
		16#1124# => X"a86b0000",
		16#1125# => X"04000633",
		16#1126# => X"a842758c",
		16#1127# => X"18600001",
		16#1128# => X"d401581c",
		16#1129# => X"d4016020",
		16#112a# => X"04001124",
		16#112b# => X"a8633cef",
		16#112c# => X"18800001",
		16#112d# => X"846200a8",
		16#112e# => X"a884758c",
		16#112f# => X"844200a0",
		16#1130# => X"84a400a4",
		16#1131# => X"18800001",
		16#1132# => X"d4011004",
		16#1133# => X"a8843c34",
		16#1134# => X"d4012808",
		16#1135# => X"04000623",
		16#1136# => X"d4012000",
		16#1137# => X"18a00001",
		16#1138# => X"a8620000",
		16#1139# => X"a8a5758c",
		16#113a# => X"848500ac",
		16#113b# => X"844500b0",
		16#113c# => X"d401580c",
		16#113d# => X"d4016010",
		16#113e# => X"d4012014",
		16#113f# => X"0400058c",
		16#1140# => X"d4011018",
		16#1141# => X"847200a0",
		16#1142# => X"04000589",
		16#1143# => X"a84b0000",
		16#1144# => X"a8620000",
		16#1145# => X"040003db",
		16#1146# => X"a88b0000",
		16#1147# => X"04000611",
		16#1148# => X"a86b0000",
		16#1149# => X"18600001",
		16#114a# => X"d401581c",
		16#114b# => X"d4016020",
		16#114c# => X"04001102",
		16#114d# => X"a8633cef",
		16#114e# => X"18800001",
		16#114f# => X"847e00a8",
		16#1150# => X"84be00a4",
		16#1151# => X"845e00a0",
		16#1152# => X"a8843c3b",
		16#1153# => X"d4012808",
		16#1154# => X"d4011004",
		16#1155# => X"04000603",
		16#1156# => X"d4012000",
		16#1157# => X"849e00ac",
		16#1158# => X"a8620000",
		16#1159# => X"845e00b0",
		16#115a# => X"d401580c",
		16#115b# => X"d4016010",
		16#115c# => X"d4012014",
		16#115d# => X"0400056e",
		16#115e# => X"d4011018",
		16#115f# => X"847000a0",
		16#1160# => X"0400056b",
		16#1161# => X"a84b0000",
		16#1162# => X"a8620000",
		16#1163# => X"040003bd",
		16#1164# => X"a88b0000",
		16#1165# => X"040005f3",
		16#1166# => X"a86b0000",
		16#1167# => X"18600001",
		16#1168# => X"d401581c",
		16#1169# => X"d4016020",
		16#116a# => X"040010e4",
		16#116b# => X"a8633cef",
		16#116c# => X"18800001",
		16#116d# => X"847c00a8",
		16#116e# => X"84bc00a4",
		16#116f# => X"845c00a0",
		16#1170# => X"a8843c42",
		16#1171# => X"d4012808",
		16#1172# => X"d4011004",
		16#1173# => X"040005e5",
		16#1174# => X"d4012000",
		16#1175# => X"849c00ac",
		16#1176# => X"a8620000",
		16#1177# => X"845c00b0",
		16#1178# => X"d401580c",
		16#1179# => X"d4016010",
		16#117a# => X"d4012014",
		16#117b# => X"04000550",
		16#117c# => X"d4011018",
		16#117d# => X"847000a0",
		16#117e# => X"0400054d",
		16#117f# => X"a84b0000",
		16#1180# => X"a8620000",
		16#1181# => X"0400039f",
		16#1182# => X"a88b0000",
		16#1183# => X"040005d5",
		16#1184# => X"a86b0000",
		16#1185# => X"18600001",
		16#1186# => X"d401581c",
		16#1187# => X"d4016020",
		16#1188# => X"040010c6",
		16#1189# => X"a8633cef",
		16#118a# => X"18800001",
		16#118b# => X"847a00a8",
		16#118c# => X"84ba00a4",
		16#118d# => X"845a00a0",
		16#118e# => X"a8843c49",
		16#118f# => X"d4012808",
		16#1190# => X"d4011004",
		16#1191# => X"040005c7",
		16#1192# => X"d4012000",
		16#1193# => X"849a00ac",
		16#1194# => X"a8620000",
		16#1195# => X"845a00b0",
		16#1196# => X"d401580c",
		16#1197# => X"d4016010",
		16#1198# => X"d4012014",
		16#1199# => X"04000532",
		16#119a# => X"d4011018",
		16#119b# => X"846e00a0",
		16#119c# => X"0400052f",
		16#119d# => X"a84b0000",
		16#119e# => X"a8620000",
		16#119f# => X"04000381",
		16#11a0# => X"a88b0000",
		16#11a1# => X"040005b7",
		16#11a2# => X"a86b0000",
		16#11a3# => X"18600001",
		16#11a4# => X"d401581c",
		16#11a5# => X"d4016020",
		16#11a6# => X"040010a8",
		16#11a7# => X"a8633cef",
		16#11a8# => X"18800001",
		16#11a9# => X"847800a8",
		16#11aa# => X"84b800a4",
		16#11ab# => X"845800a0",
		16#11ac# => X"a8843c50",
		16#11ad# => X"d4012808",
		16#11ae# => X"d4011004",
		16#11af# => X"040005a9",
		16#11b0# => X"d4012000",
		16#11b1# => X"849800ac",
		16#11b2# => X"a8620000",
		16#11b3# => X"845800b0",
		16#11b4# => X"d401580c",
		16#11b5# => X"d4016010",
		16#11b6# => X"d4012014",
		16#11b7# => X"04000514",
		16#11b8# => X"d4011018",
		16#11b9# => X"846e00a0",
		16#11ba# => X"04000511",
		16#11bb# => X"a84b0000",
		16#11bc# => X"a8620000",
		16#11bd# => X"04000363",
		16#11be# => X"a88b0000",
		16#11bf# => X"04000599",
		16#11c0# => X"a86b0000",
		16#11c1# => X"18600001",
		16#11c2# => X"d401581c",
		16#11c3# => X"d4016020",
		16#11c4# => X"0400108a",
		16#11c5# => X"a8633cef",
		16#11c6# => X"84560000",
		16#11c7# => X"84760008",
		16#11c8# => X"84960004",
		16#11c9# => X"d4011004",
		16#11ca# => X"18400001",
		16#11cb# => X"d4012008",
		16#11cc# => X"a8423d3b",
		16#11cd# => X"0400058b",
		16#11ce# => X"d4011000",
		16#11cf# => X"18600001",
		16#11d0# => X"8496000c",
		16#11d1# => X"84560010",
		16#11d2# => X"a8633d18",
		16#11d3# => X"d401580c",
		16#11d4# => X"d4016010",
		16#11d5# => X"d4012014",
		16#11d6# => X"04001078",
		16#11d7# => X"d4011018",
		16#11d8# => X"18400001",
		16#11d9# => X"84740008",
		16#11da# => X"84940004",
		16#11db# => X"84b40000",
		16#11dc# => X"a8423d3f",
		16#11dd# => X"d4012804",
		16#11de# => X"d4011000",
		16#11df# => X"04000579",
		16#11e0# => X"d4012008",
		16#11e1# => X"18600001",
		16#11e2# => X"84540010",
		16#11e3# => X"8494000c",
		16#11e4# => X"a8633d18",
		16#11e5# => X"d4011018",
		16#11e6# => X"d401580c",
		16#11e7# => X"d4016010",
		16#11e8# => X"04001066",
		16#11e9# => X"d4012014",
		16#11ea# => X"9c210054",
		16#11eb# => X"8521fffc",
		16#11ec# => X"8441ffd4",
		16#11ed# => X"85c1ffd8",
		16#11ee# => X"8601ffdc",
		16#11ef# => X"8641ffe0",
		16#11f0# => X"8681ffe4",
		16#11f1# => X"86c1ffe8",
		16#11f2# => X"8701ffec",
		16#11f3# => X"8741fff0",
		16#11f4# => X"8781fff4",
		16#11f5# => X"44004800",
		16#11f6# => X"87c1fff8",
		16#11f7# => X"d7e177ec",
		16#11f8# => X"d7e187f0",
		16#11f9# => X"d7e197f4",
		16#11fa# => X"d7e14ffc",
		16#11fb# => X"d7e117e8",
		16#11fc# => X"d7e1a7f8",
		16#11fd# => X"a9c40000",
		16#11fe# => X"9c21ffd8",
		16#11ff# => X"aa030000",
		16#1200# => X"bda40000",
		16#1201# => X"10000012",
		16#1202# => X"aa460000",
		16#1203# => X"a860c7ff",
		16#1204# => X"9c400000",
		16#1205# => X"e2851800",
		16#1206# => X"9c420001",
		16#1207# => X"04000fe4",
		16#1208# => X"e0741000",
		16#1209# => X"18600001",
		16#120a# => X"d4018000",
		16#120b# => X"a8633d44",
		16#120c# => X"d4019004",
		16#120d# => X"d4011008",
		16#120e# => X"04001040",
		16#120f# => X"d401580c",
		16#1210# => X"e54e1000",
		16#1211# => X"13fffff6",
		16#1212# => X"9c420001",
		16#1213# => X"9c210028",
		16#1214# => X"8521fffc",
		16#1215# => X"8441ffe8",
		16#1216# => X"85c1ffec",
		16#1217# => X"8601fff0",
		16#1218# => X"8641fff4",
		16#1219# => X"44004800",
		16#121a# => X"8681fff8",
		16#121b# => X"d7e117f0",
		16#121c# => X"d7e177f4",
		16#121d# => X"d7e187f8",
		16#121e# => X"d7e14ffc",
		16#121f# => X"1a000001",
		16#1220# => X"9c21ffe0",
		16#1221# => X"07fff7f9",
		16#1222# => X"9dc00000",
		16#1223# => X"aa103d63",
		16#1224# => X"a84b0000",
		16#1225# => X"a880c8ff",
		16#1226# => X"9dce0001",
		16#1227# => X"04000fc4",
		16#1228# => X"e06e2000",
		16#1229# => X"18600001",
		16#122a# => X"d4011000",
		16#122b# => X"a8633d44",
		16#122c# => X"d4018004",
		16#122d# => X"d4017008",
		16#122e# => X"04001020",
		16#122f# => X"d401580c",
		16#1230# => X"bc2e0020",
		16#1231# => X"13fffff5",
		16#1232# => X"a880c8ff",
		16#1233# => X"1a000001",
		16#1234# => X"9dc00000",
		16#1235# => X"aa103d6d",
		16#1236# => X"a880c93f",
		16#1237# => X"9dce0001",
		16#1238# => X"04000fb3",
		16#1239# => X"e06e2000",
		16#123a# => X"18600001",
		16#123b# => X"d4011000",
		16#123c# => X"a8633d44",
		16#123d# => X"d4018004",
		16#123e# => X"d4017008",
		16#123f# => X"0400100f",
		16#1240# => X"d401580c",
		16#1241# => X"bc2e0020",
		16#1242# => X"13fffff5",
		16#1243# => X"a880c93f",
		16#1244# => X"1a000001",
		16#1245# => X"9dc00000",
		16#1246# => X"aa103c30",
		16#1247# => X"a880c9ff",
		16#1248# => X"9dce0001",
		16#1249# => X"04000fa2",
		16#124a# => X"e06e2000",
		16#124b# => X"18600001",
		16#124c# => X"d4011000",
		16#124d# => X"a8633d44",
		16#124e# => X"d4018004",
		16#124f# => X"d4017008",
		16#1250# => X"04000ffe",
		16#1251# => X"d401580c",
		16#1252# => X"bc2e0020",
		16#1253# => X"13fffff5",
		16#1254# => X"a880c9ff",
		16#1255# => X"1a000001",
		16#1256# => X"9dc00000",
		16#1257# => X"aa103c2d",
		16#1258# => X"a880cabf",
		16#1259# => X"9dce0001",
		16#125a# => X"04000f91",
		16#125b# => X"e06e2000",
		16#125c# => X"18600001",
		16#125d# => X"d4011000",
		16#125e# => X"a8633d44",
		16#125f# => X"d4018004",
		16#1260# => X"d4017008",
		16#1261# => X"04000fed",
		16#1262# => X"d401580c",
		16#1263# => X"bc2e0020",
		16#1264# => X"13fffff5",
		16#1265# => X"a880cabf",
		16#1266# => X"1a000001",
		16#1267# => X"9dc00000",
		16#1268# => X"aa103c34",
		16#1269# => X"a880caff",
		16#126a# => X"9dce0001",
		16#126b# => X"04000f80",
		16#126c# => X"e06e2000",
		16#126d# => X"18600001",
		16#126e# => X"d4011000",
		16#126f# => X"a8633d44",
		16#1270# => X"d4018004",
		16#1271# => X"d4017008",
		16#1272# => X"04000fdc",
		16#1273# => X"d401580c",
		16#1274# => X"bc2e0020",
		16#1275# => X"13fffff5",
		16#1276# => X"a880caff",
		16#1277# => X"1a000001",
		16#1278# => X"9dc00000",
		16#1279# => X"aa103c3b",
		16#127a# => X"a880cb3f",
		16#127b# => X"9dce0001",
		16#127c# => X"04000f6f",
		16#127d# => X"e06e2000",
		16#127e# => X"18600001",
		16#127f# => X"d4011000",
		16#1280# => X"a8633d44",
		16#1281# => X"d4018004",
		16#1282# => X"d4017008",
		16#1283# => X"04000fcb",
		16#1284# => X"d401580c",
		16#1285# => X"bc2e0020",
		16#1286# => X"13fffff5",
		16#1287# => X"a880cb3f",
		16#1288# => X"1a000001",
		16#1289# => X"9dc00000",
		16#128a# => X"aa103c42",
		16#128b# => X"a880cb7f",
		16#128c# => X"9dce0001",
		16#128d# => X"04000f5e",
		16#128e# => X"e06e2000",
		16#128f# => X"18600001",
		16#1290# => X"d4011000",
		16#1291# => X"a8633d44",
		16#1292# => X"d4018004",
		16#1293# => X"d4017008",
		16#1294# => X"04000fba",
		16#1295# => X"d401580c",
		16#1296# => X"bc2e0020",
		16#1297# => X"13fffff5",
		16#1298# => X"a880cb7f",
		16#1299# => X"1a000001",
		16#129a# => X"9dc00000",
		16#129b# => X"aa103c49",
		16#129c# => X"a880cbbf",
		16#129d# => X"9dce0001",
		16#129e# => X"04000f4d",
		16#129f# => X"e06e2000",
		16#12a0# => X"18600001",
		16#12a1# => X"d4011000",
		16#12a2# => X"a8633d44",
		16#12a3# => X"d4018004",
		16#12a4# => X"d4017008",
		16#12a5# => X"04000fa9",
		16#12a6# => X"d401580c",
		16#12a7# => X"bc2e0020",
		16#12a8# => X"13fffff5",
		16#12a9# => X"a880cbbf",
		16#12aa# => X"1a000001",
		16#12ab# => X"9dc00000",
		16#12ac# => X"aa103c50",
		16#12ad# => X"a880cbff",
		16#12ae# => X"9dce0001",
		16#12af# => X"04000f3c",
		16#12b0# => X"e06e2000",
		16#12b1# => X"18600001",
		16#12b2# => X"d4011000",
		16#12b3# => X"a8633d44",
		16#12b4# => X"d4018004",
		16#12b5# => X"d4017008",
		16#12b6# => X"04000f98",
		16#12b7# => X"d401580c",
		16#12b8# => X"bc2e0020",
		16#12b9# => X"13fffff5",
		16#12ba# => X"a880cbff",
		16#12bb# => X"9c210020",
		16#12bc# => X"8521fffc",
		16#12bd# => X"8441fff0",
		16#12be# => X"85c1fff4",
		16#12bf# => X"44004800",
		16#12c0# => X"8601fff8",
		16#12c1# => X"9c21fffc",
		16#12c2# => X"d4014800",
		16#12c3# => X"9d600000",
		16#12c4# => X"9d040000",
		16#12c5# => X"9ca30000",
		16#12c6# => X"e4285800",
		16#12c7# => X"0c000036",
		16#12c8# => X"9ce00000",
		16#12c9# => X"e4482800",
		16#12ca# => X"10000032",
		16#12cb# => X"e4082800",
		16#12cc# => X"1000002e",
		16#12cd# => X"e48b4000",
		16#12ce# => X"0c00000d",
		16#12cf# => X"9da00020",
		16#12d0# => X"19208000",
		16#12d1# => X"9cc0ffff",
		16#12d2# => X"e0654803",
		16#12d3# => X"b8870001",
		16#12d4# => X"9de50000",
		16#12d5# => X"b863005f",
		16#12d6# => X"e1ad3000",
		16#12d7# => X"e0e41804",
		16#12d8# => X"e4874000",
		16#12d9# => X"13fffff9",
		16#12da# => X"b8a50001",
		16#12db# => X"b8e70041",
		16#12dc# => X"9dad0001",
		16#12dd# => X"9d200000",
		16#12de# => X"e4896800",
		16#12df# => X"0c00001e",
		16#12e0# => X"9caf0000",
		16#12e1# => X"19e08000",
		16#12e2# => X"9e200000",
		16#12e3# => X"e0657803",
		16#12e4# => X"b8870001",
		16#12e5# => X"b863005f",
		16#12e6# => X"e0e41804",
		16#12e7# => X"e0c74002",
		16#12e8# => X"e0667803",
		16#12e9# => X"b863005f",
		16#12ea# => X"9c800000",
		16#12eb# => X"e4232000",
		16#12ec# => X"10000003",
		16#12ed# => X"b86b0001",
		16#12ee# => X"9c800001",
		16#12ef# => X"b8a50001",
		16#12f0# => X"e4248800",
		16#12f1# => X"0c000003",
		16#12f2# => X"e1632004",
		16#12f3# => X"9ce60000",
		16#12f4# => X"9d290001",
		16#12f5# => X"e4896800",
		16#12f6# => X"13ffffed",
		16#12f7# => X"15000000",
		16#12f8# => X"00000005",
		16#12f9# => X"15000000",
		16#12fa# => X"00000003",
		16#12fb# => X"9d600001",
		16#12fc# => X"9ce50000",
		16#12fd# => X"85210000",
		16#12fe# => X"44004800",
		16#12ff# => X"9c210004",
		16#1300# => X"9c21fff8",
		16#1301# => X"d4014800",
		16#1302# => X"d4017004",
		16#1303# => X"9ca30000",
		16#1304# => X"9dc00000",
		16#1305# => X"e5850000",
		16#1306# => X"0c000004",
		16#1307# => X"9c600000",
		16#1308# => X"9dc00001",
		16#1309# => X"e0a02802",
		16#130a# => X"e5840000",
		16#130b# => X"0c000004",
		16#130c# => X"15000000",
		16#130d# => X"9dce0001",
		16#130e# => X"e0802002",
		16#130f# => X"07ffffb2",
		16#1310# => X"9c650000",
		16#1311# => X"bc0e0001",
		16#1312# => X"0c000003",
		16#1313# => X"15000000",
		16#1314# => X"e1605802",
		16#1315# => X"85210000",
		16#1316# => X"85c10004",
		16#1317# => X"44004800",
		16#1318# => X"9c210008",
		16#1319# => X"d7e117fc",
		16#131a# => X"84c30000",
		16#131b# => X"bca60001",
		16#131c# => X"1000004e",
		16#131d# => X"9c21fffc",
		16#131e# => X"84e40000",
		16#131f# => X"bca70001",
		16#1320# => X"1000006e",
		16#1321# => X"bc260004",
		16#1322# => X"0c000083",
		16#1323# => X"bc070004",
		16#1324# => X"1000006a",
		16#1325# => X"bc270002",
		16#1326# => X"0c000055",
		16#1327# => X"bc060002",
		16#1328# => X"10000066",
		16#1329# => X"15000000",
		16#132a# => X"84e30008",
		16#132b# => X"85a40008",
		16#132c# => X"8583000c",
		16#132d# => X"e1676802",
		16#132e# => X"b9eb009f",
		16#132f# => X"e0cf5805",
		16#1330# => X"e0c67802",
		16#1331# => X"bd46001f",
		16#1332# => X"1000003c",
		16#1333# => X"8504000c",
		16#1334# => X"bdab0000",
		16#1335# => X"10000064",
		16#1336# => X"9da00001",
		16#1337# => X"e1683048",
		16#1338# => X"e0cd3008",
		16#1339# => X"9cc6ffff",
		16#133a# => X"e1064003",
		16#133b# => X"e0c04002",
		16#133c# => X"e1064004",
		16#133d# => X"b908005f",
		16#133e# => X"e1085804",
		16#133f# => X"84630004",
		16#1340# => X"84840004",
		16#1341# => X"e4032000",
		16#1342# => X"10000035",
		16#1343# => X"e0886000",
		16#1344# => X"bc030000",
		16#1345# => X"10000003",
		16#1346# => X"e08c4002",
		16#1347# => X"e0886002",
		16#1348# => X"bd840000",
		16#1349# => X"1000004a",
		16#134a# => X"9c400000",
		16#134b# => X"d4053808",
		16#134c# => X"d4051004",
		16#134d# => X"d405200c",
		16#134e# => X"18403fff",
		16#134f# => X"9c64ffff",
		16#1350# => X"a842fffe",
		16#1351# => X"e4431000",
		16#1352# => X"1000000d",
		16#1353# => X"9cc00003",
		16#1354# => X"84650008",
		16#1355# => X"e0842000",
		16#1356# => X"18403fff",
		16#1357# => X"9cc4ffff",
		16#1358# => X"a842fffe",
		16#1359# => X"e4a61000",
		16#135a# => X"13fffffb",
		16#135b# => X"9c63ffff",
		16#135c# => X"d405200c",
		16#135d# => X"d4051808",
		16#135e# => X"9cc00003",
		16#135f# => X"a8650000",
		16#1360# => X"bd640000",
		16#1361# => X"10000009",
		16#1362# => X"d4053000",
		16#1363# => X"b8c40041",
		16#1364# => X"84a50008",
		16#1365# => X"a4840001",
		16#1366# => X"9ca50001",
		16#1367# => X"e0843004",
		16#1368# => X"d4032808",
		16#1369# => X"d403200c",
		16#136a# => X"9c210004",
		16#136b# => X"a9630000",
		16#136c# => X"44004800",
		16#136d# => X"8441fffc",
		16#136e# => X"e5a76800",
		16#136f# => X"1000001c",
		16#1370# => X"15000000",
		16#1371# => X"84630004",
		16#1372# => X"84840004",
		16#1373# => X"e4032000",
		16#1374# => X"0fffffd0",
		16#1375# => X"9d000000",
		16#1376# => X"e0886000",
		16#1377# => X"d4051804",
		16#1378# => X"d4053808",
		16#1379# => X"03ffffe5",
		16#137a# => X"d405200c",
		16#137b# => X"bc260002",
		16#137c# => X"13ffffee",
		16#137d# => X"15000000",
		16#137e# => X"d4053000",
		16#137f# => X"84c30004",
		16#1380# => X"d4053004",
		16#1381# => X"84c30008",
		16#1382# => X"d4053008",
		16#1383# => X"84c3000c",
		16#1384# => X"d405300c",
		16#1385# => X"84c30004",
		16#1386# => X"84840004",
		16#1387# => X"a8650000",
		16#1388# => X"e0843003",
		16#1389# => X"03ffffe1",
		16#138a# => X"d4052004",
		16#138b# => X"a8ed0000",
		16#138c# => X"03ffffb3",
		16#138d# => X"9d800000",
		16#138e# => X"a8640000",
		16#138f# => X"9c210004",
		16#1390# => X"a9630000",
		16#1391# => X"44004800",
		16#1392# => X"8441fffc",
		16#1393# => X"e0802002",
		16#1394# => X"9c600001",
		16#1395# => X"d4053808",
		16#1396# => X"d4051804",
		16#1397# => X"03ffffb7",
		16#1398# => X"d405200c",
		16#1399# => X"bc0b0000",
		16#139a# => X"13ffffa5",
		16#139b# => X"e16c3048",
		16#139c# => X"e1ad3008",
		16#139d# => X"e0e73000",
		16#139e# => X"9ccdffff",
		16#139f# => X"e1866003",
		16#13a0# => X"e0c06002",
		16#13a1# => X"e1866004",
		16#13a2# => X"b98c005f",
		16#13a3# => X"03ffff9c",
		16#13a4# => X"e18c5804",
		16#13a5# => X"bc270004",
		16#13a6# => X"13ffffc4",
		16#13a7# => X"15000000",
		16#13a8# => X"84a30004",
		16#13a9# => X"84840004",
		16#13aa# => X"e4252000",
		16#13ab# => X"0fffffbf",
		16#13ac# => X"15000000",
		16#13ad# => X"18600001",
		16#13ae# => X"03ffffbc",
		16#13af# => X"a8633d7c",
		16#13b0# => X"d7e117fc",
		16#13b1# => X"84a30000",
		16#13b2# => X"9c21fffc",
		16#13b3# => X"8483000c",
		16#13b4# => X"bc450001",
		16#13b5# => X"0c00003d",
		16#13b6# => X"84c30004",
		16#13b7# => X"bc050004",
		16#13b8# => X"10000037",
		16#13b9# => X"bc050002",
		16#13ba# => X"10000024",
		16#13bb# => X"bc040000",
		16#13bc# => X"1000001b",
		16#13bd# => X"15000000",
		16#13be# => X"84630008",
		16#13bf# => X"bd63ff82",
		16#13c0# => X"0c000039",
		16#13c1# => X"bd43007f",
		16#13c2# => X"1000002d",
		16#13c3# => X"a4a4007f",
		16#13c4# => X"bc250040",
		16#13c5# => X"0c000021",
		16#13c6# => X"9c63007f",
		16#13c7# => X"9c84003f",
		16#13c8# => X"bd640000",
		16#13c9# => X"0c000023",
		16#13ca# => X"15000000",
		16#13cb# => X"1840007f",
		16#13cc# => X"b8a40047",
		16#13cd# => X"a842ffff",
		16#13ce# => X"a48300ff",
		16#13cf# => X"e0651003",
		16#13d0# => X"b8840017",
		16#13d1# => X"b8a6001f",
		16#13d2# => X"e0832004",
		16#13d3# => X"9c210004",
		16#13d4# => X"e1642804",
		16#13d5# => X"44004800",
		16#13d6# => X"8441fffc",
		16#13d7# => X"a8640000",
		16#13d8# => X"b8a6001f",
		16#13d9# => X"e0832004",
		16#13da# => X"9c210004",
		16#13db# => X"e1642804",
		16#13dc# => X"44004800",
		16#13dd# => X"8441fffc",
		16#13de# => X"9c800000",
		16#13df# => X"b8a6001f",
		16#13e0# => X"a8640000",
		16#13e1# => X"9c210004",
		16#13e2# => X"e0832004",
		16#13e3# => X"8441fffc",
		16#13e4# => X"44004800",
		16#13e5# => X"e1642804",
		16#13e6# => X"a4a40080",
		16#13e7# => X"bc050000",
		16#13e8# => X"13ffffe1",
		16#13e9# => X"bd640000",
		16#13ea# => X"03ffffde",
		16#13eb# => X"9c840040",
		16#13ec# => X"b8840041",
		16#13ed# => X"03ffffde",
		16#13ee# => X"9c630001",
		16#13ef# => X"18807f80",
		16#13f0# => X"03ffffe1",
		16#13f1# => X"9c600000",
		16#13f2# => X"18400010",
		16#13f3# => X"e0641004",
		16#13f4# => X"1840007f",
		16#13f5# => X"18807f80",
		16#13f6# => X"a842ffff",
		16#13f7# => X"03ffffda",
		16#13f8# => X"e0631003",
		16#13f9# => X"9ce0ff82",
		16#13fa# => X"e0671802",
		16#13fb# => X"bd430019",
		16#13fc# => X"1000001f",
		16#13fd# => X"9ca00000",
		16#13fe# => X"9ce00001",
		16#13ff# => X"e0a41848",
		16#1400# => X"e0671808",
		16#1401# => X"9c63ffff",
		16#1402# => X"e0832003",
		16#1403# => X"e0602002",
		16#1404# => X"e0632004",
		16#1405# => X"b863005f",
		16#1406# => X"e0a32804",
		16#1407# => X"a465007f",
		16#1408# => X"bc230040",
		16#1409# => X"10000012",
		16#140a# => X"15000000",
		16#140b# => X"a4650080",
		16#140c# => X"bc030000",
		16#140d# => X"10000004",
		16#140e# => X"18403fff",
		16#140f# => X"9ca50040",
		16#1410# => X"18403fff",
		16#1411# => X"b8650047",
		16#1412# => X"a842ffff",
		16#1413# => X"9c800001",
		16#1414# => X"e4451000",
		16#1415# => X"1840007f",
		16#1416# => X"a842ffff",
		16#1417# => X"13ffffb9",
		16#1418# => X"e0631003",
		16#1419# => X"03ffffb7",
		16#141a# => X"9c800000",
		16#141b# => X"03fffff5",
		16#141c# => X"9ca5003f",
		16#141d# => X"d7e117fc",
		16#141e# => X"1840007f",
		16#141f# => X"84a30000",
		16#1420# => X"a842ffff",
		16#1421# => X"b8c50057",
		16#1422# => X"b8e5005f",
		16#1423# => X"9c21fffc",
		16#1424# => X"a4c600ff",
		16#1425# => X"d4043804",
		16#1426# => X"bc260000",
		16#1427# => X"10000016",
		16#1428# => X"e0651003",
		16#1429# => X"bc230000",
		16#142a# => X"0c000020",
		16#142b# => X"9ca0ff82",
		16#142c# => X"b8630007",
		16#142d# => X"d4042808",
		16#142e# => X"9ca00003",
		16#142f# => X"d4042800",
		16#1430# => X"9ca0ff81",
		16#1431# => X"18403fff",
		16#1432# => X"e0631800",
		16#1433# => X"a842ffff",
		16#1434# => X"a8c50000",
		16#1435# => X"e4a31000",
		16#1436# => X"13fffffb",
		16#1437# => X"9ca5ffff",
		16#1438# => X"9c210004",
		16#1439# => X"d4043008",
		16#143a# => X"d404180c",
		16#143b# => X"44004800",
		16#143c# => X"8441fffc",
		16#143d# => X"bc2600ff",
		16#143e# => X"0c000011",
		16#143f# => X"9cc6ff81",
		16#1440# => X"b8630007",
		16#1441# => X"18404000",
		16#1442# => X"d4043008",
		16#1443# => X"e0631004",
		16#1444# => X"9ca00003",
		16#1445# => X"d4042800",
		16#1446# => X"d404180c",
		16#1447# => X"9c210004",
		16#1448# => X"44004800",
		16#1449# => X"8441fffc",
		16#144a# => X"9c600002",
		16#144b# => X"9c210004",
		16#144c# => X"d4041800",
		16#144d# => X"44004800",
		16#144e# => X"8441fffc",
		16#144f# => X"bc230000",
		16#1450# => X"0c00000a",
		16#1451# => X"15000000",
		16#1452# => X"18400010",
		16#1453# => X"e0a51003",
		16#1454# => X"bc050000",
		16#1455# => X"13fffff0",
		16#1456# => X"15000000",
		16#1457# => X"9ca00001",
		16#1458# => X"03ffffee",
		16#1459# => X"d4042800",
		16#145a# => X"9c600004",
		16#145b# => X"03ffffec",
		16#145c# => X"d4041800",
		16#145d# => X"d7e14ffc",
		16#145e# => X"d7e117f4",
		16#145f# => X"d7e177f8",
		16#1460# => X"9c21ffbc",
		16#1461# => X"9dc10020",
		16#1462# => X"d4011834",
		16#1463# => X"d4012030",
		16#1464# => X"9c610034",
		16#1465# => X"a88e0000",
		16#1466# => X"07ffffb7",
		16#1467# => X"9c410010",
		16#1468# => X"9c610030",
		16#1469# => X"07ffffb4",
		16#146a# => X"a8820000",
		16#146b# => X"a86e0000",
		16#146c# => X"a8820000",
		16#146d# => X"07fffeac",
		16#146e# => X"a8a10000",
		16#146f# => X"07ffff41",
		16#1470# => X"a86b0000",
		16#1471# => X"9c210044",
		16#1472# => X"8521fffc",
		16#1473# => X"8441fff4",
		16#1474# => X"44004800",
		16#1475# => X"85c1fff8",
		16#1476# => X"d7e14ffc",
		16#1477# => X"d7e117f4",
		16#1478# => X"d7e177f8",
		16#1479# => X"9c21ffbc",
		16#147a# => X"9dc10020",
		16#147b# => X"d4011834",
		16#147c# => X"d4012030",
		16#147d# => X"9c610034",
		16#147e# => X"a88e0000",
		16#147f# => X"07ffff9e",
		16#1480# => X"9c410010",
		16#1481# => X"9c610030",
		16#1482# => X"07ffff9b",
		16#1483# => X"a8820000",
		16#1484# => X"84c10014",
		16#1485# => X"a86e0000",
		16#1486# => X"acc60001",
		16#1487# => X"a8820000",
		16#1488# => X"a8a10000",
		16#1489# => X"07fffe90",
		16#148a# => X"d4013014",
		16#148b# => X"07ffff25",
		16#148c# => X"a86b0000",
		16#148d# => X"9c210044",
		16#148e# => X"8521fffc",
		16#148f# => X"8441fff4",
		16#1490# => X"44004800",
		16#1491# => X"85c1fff8",
		16#1492# => X"d7e14ffc",
		16#1493# => X"d7e117f4",
		16#1494# => X"d7e177f8",
		16#1495# => X"9c21ffbc",
		16#1496# => X"9c410020",
		16#1497# => X"d4011834",
		16#1498# => X"d4012030",
		16#1499# => X"9c610034",
		16#149a# => X"a8820000",
		16#149b# => X"07ffff82",
		16#149c# => X"9dc10010",
		16#149d# => X"9c610030",
		16#149e# => X"07ffff7f",
		16#149f# => X"a88e0000",
		16#14a0# => X"84a10020",
		16#14a1# => X"bc450001",
		16#14a2# => X"0c00005e",
		16#14a3# => X"84c10010",
		16#14a4# => X"bc460001",
		16#14a5# => X"0c00006d",
		16#14a6# => X"bc250004",
		16#14a7# => X"0c000055",
		16#14a8# => X"bc260004",
		16#14a9# => X"0c000065",
		16#14aa# => X"bc250002",
		16#14ab# => X"0c000055",
		16#14ac# => X"bc260002",
		16#14ad# => X"0c000065",
		16#14ae# => X"9c600000",
		16#14af# => X"8481001c",
		16#14b0# => X"a8a30000",
		16#14b1# => X"04000916",
		16#14b2# => X"84c1002c",
		16#14b3# => X"84610024",
		16#14b4# => X"84410014",
		16#14b5# => X"84810028",
		16#14b6# => X"e0431005",
		16#14b7# => X"84a10018",
		16#14b8# => X"e0601002",
		16#14b9# => X"e0852000",
		16#14ba# => X"e0431004",
		16#14bb# => X"9c640002",
		16#14bc# => X"b842005f",
		16#14bd# => X"d4011808",
		16#14be# => X"bd6b0000",
		16#14bf# => X"d4011004",
		16#14c0# => X"10000008",
		16#14c1# => X"a86b0000",
		16#14c2# => X"a44b0001",
		16#14c3# => X"bc020000",
		16#14c4# => X"0c00002a",
		16#14c5# => X"9c840003",
		16#14c6# => X"b86b0041",
		16#14c7# => X"d4012008",
		16#14c8# => X"18403fff",
		16#14c9# => X"a842ffff",
		16#14ca# => X"e4431000",
		16#14cb# => X"10000014",
		16#14cc# => X"84810008",
		16#14cd# => X"00000008",
		16#14ce# => X"e0631800",
		16#14cf# => X"18403fff",
		16#14d0# => X"a842ffff",
		16#14d1# => X"e4a31000",
		16#14d2# => X"0c00000c",
		16#14d3# => X"e18c6000",
		16#14d4# => X"e0631800",
		16#14d5# => X"bd6c0000",
		16#14d6# => X"13fffff9",
		16#14d7# => X"9c84ffff",
		16#14d8# => X"18403fff",
		16#14d9# => X"a8630001",
		16#14da# => X"a842ffff",
		16#14db# => X"e4a31000",
		16#14dc# => X"13fffff8",
		16#14dd# => X"e18c6000",
		16#14de# => X"d4012008",
		16#14df# => X"a443007f",
		16#14e0# => X"bc220040",
		16#14e1# => X"0c000011",
		16#14e2# => X"a4430080",
		16#14e3# => X"9c400003",
		16#14e4# => X"d401180c",
		16#14e5# => X"d4011000",
		16#14e6# => X"a8610000",
		16#14e7# => X"07fffec9",
		16#14e8# => X"15000000",
		16#14e9# => X"9c210044",
		16#14ea# => X"8521fffc",
		16#14eb# => X"8441fff4",
		16#14ec# => X"44004800",
		16#14ed# => X"85c1fff8",
		16#14ee# => X"b98c0041",
		16#14ef# => X"18408000",
		16#14f0# => X"03ffffd6",
		16#14f1# => X"e18c1004",
		16#14f2# => X"bc220000",
		16#14f3# => X"13fffff1",
		16#14f4# => X"9c400003",
		16#14f5# => X"bc0c0000",
		16#14f6# => X"13ffffee",
		16#14f7# => X"15000000",
		16#14f8# => X"9c630040",
		16#14f9# => X"9c40ff80",
		16#14fa# => X"03ffffe9",
		16#14fb# => X"e0631003",
		16#14fc# => X"18600001",
		16#14fd# => X"bc060002",
		16#14fe# => X"13ffffe9",
		16#14ff# => X"a8633d7c",
		16#1500# => X"84810024",
		16#1501# => X"a8620000",
		16#1502# => X"84410014",
		16#1503# => X"e0441005",
		16#1504# => X"e0801002",
		16#1505# => X"e0441004",
		16#1506# => X"b842005f",
		16#1507# => X"07fffea9",
		16#1508# => X"d4011024",
		16#1509# => X"9c210044",
		16#150a# => X"8521fffc",
		16#150b# => X"8441fff4",
		16#150c# => X"44004800",
		16#150d# => X"85c1fff8",
		16#150e# => X"18600001",
		16#150f# => X"bc050002",
		16#1510# => X"13ffffd7",
		16#1511# => X"a8633d7c",
		16#1512# => X"84410014",
		16#1513# => X"84810024",
		16#1514# => X"a86e0000",
		16#1515# => X"e0441005",
		16#1516# => X"e0801002",
		16#1517# => X"e0441004",
		16#1518# => X"b842005f",
		16#1519# => X"07fffe97",
		16#151a# => X"d4011014",
		16#151b# => X"9c210044",
		16#151c# => X"8521fffc",
		16#151d# => X"8441fff4",
		16#151e# => X"44004800",
		16#151f# => X"85c1fff8",
		16#1520# => X"d7e14ffc",
		16#1521# => X"d7e117f4",
		16#1522# => X"d7e177f8",
		16#1523# => X"9c21ffcc",
		16#1524# => X"9c410010",
		16#1525# => X"d4011824",
		16#1526# => X"d4012020",
		16#1527# => X"9c610024",
		16#1528# => X"07fffef5",
		16#1529# => X"a8820000",
		16#152a# => X"9c610020",
		16#152b# => X"07fffef2",
		16#152c# => X"a8810000",
		16#152d# => X"84a10010",
		16#152e# => X"bca50001",
		16#152f# => X"1000002c",
		16#1530# => X"a8620000",
		16#1531# => X"84c10000",
		16#1532# => X"bca60001",
		16#1533# => X"10000028",
		16#1534# => X"a8610000",
		16#1535# => X"84810014",
		16#1536# => X"84610004",
		16#1537# => X"bc050004",
		16#1538# => X"e0641805",
		16#1539# => X"1000002d",
		16#153a# => X"d4011814",
		16#153b# => X"bc250002",
		16#153c# => X"0c00002a",
		16#153d# => X"bc260004",
		16#153e# => X"0c000040",
		16#153f# => X"bc260002",
		16#1540# => X"0c000035",
		16#1541# => X"84a10018",
		16#1542# => X"84810008",
		16#1543# => X"8461001c",
		16#1544# => X"e0852002",
		16#1545# => X"84e1000c",
		16#1546# => X"e4633800",
		16#1547# => X"0c00001b",
		16#1548# => X"d4012018",
		16#1549# => X"9ca0001f",
		16#154a# => X"18c04000",
		16#154b# => X"9d000000",
		16#154c# => X"e4471800",
		16#154d# => X"10000004",
		16#154e# => X"9ca5ffff",
		16#154f# => X"e1083004",
		16#1550# => X"e0633802",
		16#1551# => X"b8c60041",
		16#1552# => X"bc250000",
		16#1553# => X"13fffff9",
		16#1554# => X"e0631800",
		16#1555# => X"a488007f",
		16#1556# => X"bc240040",
		16#1557# => X"0c000015",
		16#1558# => X"a4880080",
		16#1559# => X"d401401c",
		16#155a# => X"a8620000",
		16#155b# => X"07fffe55",
		16#155c# => X"15000000",
		16#155d# => X"9c210034",
		16#155e# => X"8521fffc",
		16#155f# => X"8441fff4",
		16#1560# => X"44004800",
		16#1561# => X"85c1fff8",
		16#1562# => X"9c84ffff",
		16#1563# => X"e0631800",
		16#1564# => X"03ffffe5",
		16#1565# => X"d4012018",
		16#1566# => X"18600001",
		16#1567# => X"e4053000",
		16#1568# => X"0ffffff2",
		16#1569# => X"a8633d7c",
		16#156a# => X"03fffff1",
		16#156b# => X"15000000",
		16#156c# => X"bc240000",
		16#156d# => X"13ffffec",
		16#156e# => X"bc030000",
		16#156f# => X"13ffffea",
		16#1570# => X"9c60ff80",
		16#1571# => X"9d080040",
		16#1572# => X"e1081803",
		16#1573# => X"03ffffe7",
		16#1574# => X"d401401c",
		16#1575# => X"a8620000",
		16#1576# => X"9c400004",
		16#1577# => X"07fffe39",
		16#1578# => X"d4011010",
		16#1579# => X"9c210034",
		16#157a# => X"8521fffc",
		16#157b# => X"8441fff4",
		16#157c# => X"44004800",
		16#157d# => X"85c1fff8",
		16#157e# => X"9c600000",
		16#157f# => X"d401181c",
		16#1580# => X"d4011818",
		16#1581# => X"03ffffda",
		16#1582# => X"a8620000",
		16#1583# => X"84a30000",
		16#1584# => X"9d600001",
		16#1585# => X"e4a55800",
		16#1586# => X"10000016",
		16#1587# => X"15000000",
		16#1588# => X"84c40000",
		16#1589# => X"e4a65800",
		16#158a# => X"10000012",
		16#158b# => X"bc250004",
		16#158c# => X"0c000037",
		16#158d# => X"bc260004",
		16#158e# => X"0c000019",
		16#158f# => X"bc250002",
		16#1590# => X"0c000014",
		16#1591# => X"bc260002",
		16#1592# => X"0c00000c",
		16#1593# => X"15000000",
		16#1594# => X"84a30004",
		16#1595# => X"84c40004",
		16#1596# => X"e4053000",
		16#1597# => X"10000016",
		16#1598# => X"15000000",
		16#1599# => X"bc050000",
		16#159a# => X"0c000008",
		16#159b# => X"15000000",
		16#159c# => X"44004800",
		16#159d# => X"15000000",
		16#159e# => X"84630004",
		16#159f# => X"bc030000",
		16#15a0# => X"13fffffc",
		16#15a1# => X"15000000",
		16#15a2# => X"44004800",
		16#15a3# => X"9d60ffff",
		16#15a4# => X"bc060002",
		16#15a5# => X"13fffff7",
		16#15a6# => X"9d600000",
		16#15a7# => X"84640004",
		16#15a8# => X"bc030000",
		16#15a9# => X"13fffff3",
		16#15aa# => X"9d60ffff",
		16#15ab# => X"44004800",
		16#15ac# => X"9d600001",
		16#15ad# => X"84e30008",
		16#15ae# => X"84c40008",
		16#15af# => X"e5a73000",
		16#15b0# => X"0fffffea",
		16#15b1# => X"bc050000",
		16#15b2# => X"e5673000",
		16#15b3# => X"0c00000c",
		16#15b4# => X"bc050000",
		16#15b5# => X"84c3000c",
		16#15b6# => X"8464000c",
		16#15b7# => X"e4a61800",
		16#15b8# => X"10000004",
		16#15b9# => X"e4661800",
		16#15ba# => X"03ffffdf",
		16#15bb# => X"9d600001",
		16#15bc# => X"13ffffe0",
		16#15bd# => X"9d600000",
		16#15be# => X"bc050000",
		16#15bf# => X"0fffffec",
		16#15c0# => X"9d60ffff",
		16#15c1# => X"44004800",
		16#15c2# => X"15000000",
		16#15c3# => X"13ffffdb",
		16#15c4# => X"15000000",
		16#15c5# => X"85640004",
		16#15c6# => X"84630004",
		16#15c7# => X"44004800",
		16#15c8# => X"e16b1802",
		16#15c9# => X"d7e14ffc",
		16#15ca# => X"d7e117f4",
		16#15cb# => X"d7e177f8",
		16#15cc# => X"9c21ffcc",
		16#15cd# => X"9dc10010",
		16#15ce# => X"d4011824",
		16#15cf# => X"d4012020",
		16#15d0# => X"9c610024",
		16#15d1# => X"07fffe4c",
		16#15d2# => X"a88e0000",
		16#15d3# => X"9c610020",
		16#15d4# => X"07fffe49",
		16#15d5# => X"a8810000",
		16#15d6# => X"a86e0000",
		16#15d7# => X"07ffffac",
		16#15d8# => X"a8810000",
		16#15d9# => X"9c210034",
		16#15da# => X"8521fffc",
		16#15db# => X"8441fff4",
		16#15dc# => X"44004800",
		16#15dd# => X"85c1fff8",
		16#15de# => X"d7e14ffc",
		16#15df# => X"d7e177f8",
		16#15e0# => X"d7e117f4",
		16#15e1# => X"9c21ffcc",
		16#15e2# => X"9dc10010",
		16#15e3# => X"d4011824",
		16#15e4# => X"d4012020",
		16#15e5# => X"9c610024",
		16#15e6# => X"07fffe37",
		16#15e7# => X"a88e0000",
		16#15e8# => X"9c610020",
		16#15e9# => X"07fffe34",
		16#15ea# => X"a8810000",
		16#15eb# => X"9d600001",
		16#15ec# => X"84610010",
		16#15ed# => X"e4a35800",
		16#15ee# => X"10000007",
		16#15ef# => X"84610000",
		16#15f0# => X"e4a35800",
		16#15f1# => X"10000004",
		16#15f2# => X"a86e0000",
		16#15f3# => X"07ffff90",
		16#15f4# => X"a8810000",
		16#15f5# => X"9c210034",
		16#15f6# => X"8521fffc",
		16#15f7# => X"8441fff4",
		16#15f8# => X"44004800",
		16#15f9# => X"85c1fff8",
		16#15fa# => X"d7e14ffc",
		16#15fb# => X"d7e177f8",
		16#15fc# => X"d7e117f4",
		16#15fd# => X"9c21ffcc",
		16#15fe# => X"9dc10010",
		16#15ff# => X"d4011824",
		16#1600# => X"d4012020",
		16#1601# => X"9c610024",
		16#1602# => X"07fffe1b",
		16#1603# => X"a88e0000",
		16#1604# => X"9c610020",
		16#1605# => X"07fffe18",
		16#1606# => X"a8810000",
		16#1607# => X"9d600001",
		16#1608# => X"84610010",
		16#1609# => X"e4a35800",
		16#160a# => X"10000007",
		16#160b# => X"84610000",
		16#160c# => X"e4a35800",
		16#160d# => X"10000004",
		16#160e# => X"a86e0000",
		16#160f# => X"07ffff74",
		16#1610# => X"a8810000",
		16#1611# => X"9c210034",
		16#1612# => X"8521fffc",
		16#1613# => X"8441fff4",
		16#1614# => X"44004800",
		16#1615# => X"85c1fff8",
		16#1616# => X"d7e14ffc",
		16#1617# => X"d7e177f8",
		16#1618# => X"d7e117f4",
		16#1619# => X"9c21ffcc",
		16#161a# => X"9dc10010",
		16#161b# => X"d4011824",
		16#161c# => X"d4012020",
		16#161d# => X"9c610024",
		16#161e# => X"07fffdff",
		16#161f# => X"a88e0000",
		16#1620# => X"9c610020",
		16#1621# => X"07fffdfc",
		16#1622# => X"a8810000",
		16#1623# => X"84610010",
		16#1624# => X"bca30001",
		16#1625# => X"10000008",
		16#1626# => X"9d60ffff",
		16#1627# => X"84610000",
		16#1628# => X"bca30001",
		16#1629# => X"10000004",
		16#162a# => X"a86e0000",
		16#162b# => X"07ffff58",
		16#162c# => X"a8810000",
		16#162d# => X"9c210034",
		16#162e# => X"8521fffc",
		16#162f# => X"8441fff4",
		16#1630# => X"44004800",
		16#1631# => X"85c1fff8",
		16#1632# => X"d7e14ffc",
		16#1633# => X"d7e177f8",
		16#1634# => X"d7e117f4",
		16#1635# => X"9c21ffcc",
		16#1636# => X"9dc10010",
		16#1637# => X"d4011824",
		16#1638# => X"d4012020",
		16#1639# => X"9c610024",
		16#163a# => X"07fffde3",
		16#163b# => X"a88e0000",
		16#163c# => X"9c610020",
		16#163d# => X"07fffde0",
		16#163e# => X"a8810000",
		16#163f# => X"84610010",
		16#1640# => X"bca30001",
		16#1641# => X"10000008",
		16#1642# => X"9d60ffff",
		16#1643# => X"84610000",
		16#1644# => X"bca30001",
		16#1645# => X"10000004",
		16#1646# => X"a86e0000",
		16#1647# => X"07ffff3c",
		16#1648# => X"a8810000",
		16#1649# => X"9c210034",
		16#164a# => X"8521fffc",
		16#164b# => X"8441fff4",
		16#164c# => X"44004800",
		16#164d# => X"85c1fff8",
		16#164e# => X"d7e14ffc",
		16#164f# => X"d7e177f8",
		16#1650# => X"d7e117f4",
		16#1651# => X"9c21ffcc",
		16#1652# => X"9dc10010",
		16#1653# => X"d4011824",
		16#1654# => X"d4012020",
		16#1655# => X"9c610024",
		16#1656# => X"07fffdc7",
		16#1657# => X"a88e0000",
		16#1658# => X"9c610020",
		16#1659# => X"07fffdc4",
		16#165a# => X"a8810000",
		16#165b# => X"9d600001",
		16#165c# => X"84610010",
		16#165d# => X"e4a35800",
		16#165e# => X"10000007",
		16#165f# => X"84610000",
		16#1660# => X"e4a35800",
		16#1661# => X"10000004",
		16#1662# => X"a86e0000",
		16#1663# => X"07ffff20",
		16#1664# => X"a8810000",
		16#1665# => X"9c210034",
		16#1666# => X"8521fffc",
		16#1667# => X"8441fff4",
		16#1668# => X"44004800",
		16#1669# => X"85c1fff8",
		16#166a# => X"d7e14ffc",
		16#166b# => X"d7e177f8",
		16#166c# => X"d7e117f4",
		16#166d# => X"9c21ffcc",
		16#166e# => X"9dc10010",
		16#166f# => X"d4011824",
		16#1670# => X"d4012020",
		16#1671# => X"9c610024",
		16#1672# => X"07fffdab",
		16#1673# => X"a88e0000",
		16#1674# => X"9c610020",
		16#1675# => X"07fffda8",
		16#1676# => X"a8810000",
		16#1677# => X"9d600001",
		16#1678# => X"84610010",
		16#1679# => X"e4a35800",
		16#167a# => X"10000007",
		16#167b# => X"84610000",
		16#167c# => X"e4a35800",
		16#167d# => X"10000004",
		16#167e# => X"a86e0000",
		16#167f# => X"07ffff04",
		16#1680# => X"a8810000",
		16#1681# => X"9c210034",
		16#1682# => X"8521fffc",
		16#1683# => X"8441fff4",
		16#1684# => X"44004800",
		16#1685# => X"85c1fff8",
		16#1686# => X"d7e14ffc",
		16#1687# => X"9c21ffd4",
		16#1688# => X"d4011824",
		16#1689# => X"d4012020",
		16#168a# => X"9c610024",
		16#168b# => X"07fffd92",
		16#168c# => X"9c810010",
		16#168d# => X"9c610020",
		16#168e# => X"07fffd8f",
		16#168f# => X"a8810000",
		16#1690# => X"9d600001",
		16#1691# => X"84610010",
		16#1692# => X"e4a35800",
		16#1693# => X"10000005",
		16#1694# => X"84610000",
		16#1695# => X"e4a35800",
		16#1696# => X"0c000006",
		16#1697# => X"15000000",
		16#1698# => X"9c21002c",
		16#1699# => X"8521fffc",
		16#169a# => X"44004800",
		16#169b# => X"15000000",
		16#169c# => X"9c21002c",
		16#169d# => X"8521fffc",
		16#169e# => X"44004800",
		16#169f# => X"9d600000",
		16#16a0# => X"b883005f",
		16#16a1# => X"d7e117f8",
		16#16a2# => X"d7e14ffc",
		16#16a3# => X"9c400003",
		16#16a4# => X"9c21ffe8",
		16#16a5# => X"bc230000",
		16#16a6# => X"d4011000",
		16#16a7# => X"1000000a",
		16#16a8# => X"d4012004",
		16#16a9# => X"9c400002",
		16#16aa# => X"d4011000",
		16#16ab# => X"07fffd05",
		16#16ac# => X"a8610000",
		16#16ad# => X"9c210018",
		16#16ae# => X"8521fffc",
		16#16af# => X"44004800",
		16#16b0# => X"8441fff8",
		16#16b1# => X"a8430000",
		16#16b2# => X"9c60001e",
		16#16b3# => X"bc040000",
		16#16b4# => X"10000007",
		16#16b5# => X"d4011808",
		16#16b6# => X"18608000",
		16#16b7# => X"e4021800",
		16#16b8# => X"1000000f",
		16#16b9# => X"15000000",
		16#16ba# => X"e0401002",
		16#16bb# => X"a8620000",
		16#16bc# => X"04000750",
		16#16bd# => X"d401100c",
		16#16be# => X"9d6bffff",
		16#16bf# => X"bdab0000",
		16#16c0# => X"13ffffeb",
		16#16c1# => X"9c60001e",
		16#16c2# => X"e0425808",
		16#16c3# => X"e1635802",
		16#16c4# => X"d401100c",
		16#16c5# => X"03ffffe6",
		16#16c6# => X"d4015808",
		16#16c7# => X"18400001",
		16#16c8# => X"a8423d78",
		16#16c9# => X"03ffffe4",
		16#16ca# => X"85620000",
		16#16cb# => X"d7e117f4",
		16#16cc# => X"9c800000",
		16#16cd# => X"d7e14ffc",
		16#16ce# => X"d7e177f8",
		16#16cf# => X"9c21ffe4",
		16#16d0# => X"a8430000",
		16#16d1# => X"e4232000",
		16#16d2# => X"0c000018",
		16#16d3# => X"d4012004",
		16#16d4# => X"9c800003",
		16#16d5# => X"9dc0001e",
		16#16d6# => X"d4012000",
		16#16d7# => X"d4017008",
		16#16d8# => X"04000734",
		16#16d9# => X"d401180c",
		16#16da# => X"9d6bffff",
		16#16db# => X"bd6b0000",
		16#16dc# => X"0c000017",
		16#16dd# => X"bc0b0000",
		16#16de# => X"10000005",
		16#16df# => X"e0425808",
		16#16e0# => X"e16e5802",
		16#16e1# => X"d401100c",
		16#16e2# => X"d4015808",
		16#16e3# => X"07fffccd",
		16#16e4# => X"a8610000",
		16#16e5# => X"9c21001c",
		16#16e6# => X"8521fffc",
		16#16e7# => X"8441fff4",
		16#16e8# => X"44004800",
		16#16e9# => X"85c1fff8",
		16#16ea# => X"9c400002",
		16#16eb# => X"a8610000",
		16#16ec# => X"07fffcc4",
		16#16ed# => X"d4011000",
		16#16ee# => X"9c21001c",
		16#16ef# => X"8521fffc",
		16#16f0# => X"8441fff4",
		16#16f1# => X"44004800",
		16#16f2# => X"85c1fff8",
		16#16f3# => X"e0605802",
		16#16f4# => X"9ca00001",
		16#16f5# => X"e0821848",
		16#16f6# => X"e0651808",
		16#16f7# => X"e16e5802",
		16#16f8# => X"9c63ffff",
		16#16f9# => X"d4015808",
		16#16fa# => X"e0431003",
		16#16fb# => X"e0601002",
		16#16fc# => X"e0431004",
		16#16fd# => X"a8610000",
		16#16fe# => X"b842005f",
		16#16ff# => X"e0422004",
		16#1700# => X"07fffcb0",
		16#1701# => X"d401100c",
		16#1702# => X"9c21001c",
		16#1703# => X"8521fffc",
		16#1704# => X"8441fff4",
		16#1705# => X"44004800",
		16#1706# => X"85c1fff8",
		16#1707# => X"d7e14ffc",
		16#1708# => X"9c21ffe8",
		16#1709# => X"d4011810",
		16#170a# => X"a8810000",
		16#170b# => X"07fffd12",
		16#170c# => X"9c610010",
		16#170d# => X"84610000",
		16#170e# => X"bc030002",
		16#170f# => X"10000012",
		16#1710# => X"9d600000",
		16#1711# => X"bca30001",
		16#1712# => X"1000000f",
		16#1713# => X"bc230004",
		16#1714# => X"0c00001d",
		16#1715# => X"84610008",
		16#1716# => X"bd830000",
		16#1717# => X"1000000a",
		16#1718# => X"bda3001e",
		16#1719# => X"1000000c",
		16#171a# => X"15000000",
		16#171b# => X"84610004",
		16#171c# => X"bc030000",
		16#171d# => X"0c000018",
		16#171e# => X"15000000",
		16#171f# => X"19607fff",
		16#1720# => X"a96bffff",
		16#1721# => X"9c210018",
		16#1722# => X"8521fffc",
		16#1723# => X"44004800",
		16#1724# => X"15000000",
		16#1725# => X"9d60001e",
		16#1726# => X"e06b1802",
		16#1727# => X"8561000c",
		16#1728# => X"e16b1848",
		16#1729# => X"84610004",
		16#172a# => X"bc030000",
		16#172b# => X"13fffff6",
		16#172c# => X"15000000",
		16#172d# => X"9c210018",
		16#172e# => X"8521fffc",
		16#172f# => X"44004800",
		16#1730# => X"e1605802",
		16#1731# => X"84610004",
		16#1732# => X"e4035800",
		16#1733# => X"13ffffec",
		16#1734# => X"15000000",
		16#1735# => X"9c210018",
		16#1736# => X"8521fffc",
		16#1737# => X"44004800",
		16#1738# => X"19608000",
		16#1739# => X"d7e14ffc",
		16#173a# => X"d7e117f8",
		16#173b# => X"9c21ffe4",
		16#173c# => X"d4011810",
		16#173d# => X"a8810000",
		16#173e# => X"07fffcdf",
		16#173f# => X"9c610010",
		16#1740# => X"84810004",
		16#1741# => X"a8610000",
		16#1742# => X"e0402002",
		16#1743# => X"e0422004",
		16#1744# => X"ac42ffff",
		16#1745# => X"b842005f",
		16#1746# => X"07fffc6a",
		16#1747# => X"d4011004",
		16#1748# => X"9c21001c",
		16#1749# => X"8521fffc",
		16#174a# => X"44004800",
		16#174b# => X"8441fff8",
		16#174c# => X"d7e14ffc",
		16#174d# => X"9c21ffec",
		16#174e# => X"d4011800",
		16#174f# => X"a8610000",
		16#1750# => X"d4012004",
		16#1751# => X"d4012808",
		16#1752# => X"07fffc5e",
		16#1753# => X"d401300c",
		16#1754# => X"9c210014",
		16#1755# => X"8521fffc",
		16#1756# => X"44004800",
		16#1757# => X"15000000",
		16#1758# => X"d7e14ffc",
		16#1759# => X"d7e117f8",
		16#175a# => X"9c21ffe4",
		16#175b# => X"d4011810",
		16#175c# => X"a8810000",
		16#175d# => X"07fffcc0",
		16#175e# => X"9c610010",
		16#175f# => X"84e1000c",
		16#1760# => X"84610000",
		16#1761# => X"b8c70042",
		16#1762# => X"b8e7001e",
		16#1763# => X"84810004",
		16#1764# => X"04000636",
		16#1765# => X"84a10008",
		16#1766# => X"9c21001c",
		16#1767# => X"a84b0000",
		16#1768# => X"a86c0000",
		16#1769# => X"8521fffc",
		16#176a# => X"e1620004",
		16#176b# => X"e1830004",
		16#176c# => X"44004800",
		16#176d# => X"8441fff8",
		16#176e# => X"d7e117f8",
		16#176f# => X"d7e177fc",
		16#1770# => X"84430000",
		16#1771# => X"9c21fff8",
		16#1772# => X"bca20001",
		16#1773# => X"1000008c",
		16#1774# => X"a9630000",
		16#1775# => X"84640000",
		16#1776# => X"bca30001",
		16#1777# => X"100000cf",
		16#1778# => X"bc220004",
		16#1779# => X"0c000109",
		16#177a# => X"bc030004",
		16#177b# => X"100000cb",
		16#177c# => X"bc230002",
		16#177d# => X"0c00009a",
		16#177e# => X"bc020002",
		16#177f# => X"100000c7",
		16#1780# => X"15000000",
		16#1781# => X"858b0008",
		16#1782# => X"85e40008",
		16#1783# => X"84cb000c",
		16#1784# => X"84eb0010",
		16#1785# => X"e1ac7802",
		16#1786# => X"8444000c",
		16#1787# => X"84640010",
		16#1788# => X"ba2d009f",
		16#1789# => X"e1116805",
		16#178a# => X"e1088802",
		16#178b# => X"bd48003f",
		16#178c# => X"10000077",
		16#178d# => X"e5ac7800",
		16#178e# => X"bdad0000",
		16#178f# => X"100000bc",
		16#1790# => X"bc0d0000",
		16#1791# => X"9da8ffe0",
		16#1792# => X"bd8d0000",
		16#1793# => X"100000d4",
		16#1794# => X"a9c20000",
		16#1795# => X"9ea00000",
		16#1796# => X"e1ee6848",
		16#1797# => X"bd8d0000",
		16#1798# => X"100000dc",
		16#1799# => X"9e200001",
		16#179a# => X"9d000000",
		16#179b# => X"e1b16808",
		16#179c# => X"9e28ffff",
		16#179d# => X"e4914000",
		16#179e# => X"10000003",
		16#179f# => X"9e600001",
		16#17a0# => X"9e600000",
		16#17a1# => X"9d0dffff",
		16#17a2# => X"e2311803",
		16#17a3# => X"e1134000",
		16#17a4# => X"e1081003",
		16#17a5# => X"a8550000",
		16#17a6# => X"e1088804",
		16#17a7# => X"e1a04002",
		16#17a8# => X"e10d4004",
		16#17a9# => X"b908005f",
		16#17aa# => X"e1e87804",
		16#17ab# => X"a86f0000",
		16#17ac# => X"850b0004",
		16#17ad# => X"84840004",
		16#17ae# => X"e4082000",
		16#17af# => X"1000005d",
		16#17b0# => X"e0833800",
		16#17b1# => X"bc080000",
		16#17b2# => X"1000007f",
		16#17b3# => X"e0871802",
		16#17b4# => X"e0833802",
		16#17b5# => X"e4441800",
		16#17b6# => X"10000003",
		16#17b7# => X"9d000001",
		16#17b8# => X"9d000000",
		16#17b9# => X"e0623002",
		16#17ba# => X"e0634002",
		16#17bb# => X"bd830000",
		16#17bc# => X"1000007f",
		16#17bd# => X"9c400001",
		16#17be# => X"9d600000",
		16#17bf# => X"d4056008",
		16#17c0# => X"d4055804",
		16#17c1# => X"d405180c",
		16#17c2# => X"d4052010",
		16#17c3# => X"9cc4ffff",
		16#17c4# => X"e4862000",
		16#17c5# => X"10000003",
		16#17c6# => X"9c400001",
		16#17c7# => X"9c400000",
		16#17c8# => X"9ce3ffff",
		16#17c9# => X"19a00fff",
		16#17ca# => X"e0423800",
		16#17cb# => X"a9adffff",
		16#17cc# => X"e4426800",
		16#17cd# => X"10000020",
		16#17ce# => X"e4226800",
		16#17cf# => X"0c0000a1",
		16#17d0# => X"bc46fffe",
		16#17d1# => X"00000004",
		16#17d2# => X"84450008",
		16#17d3# => X"0c00005a",
		16#17d4# => X"bc4bfffe",
		16#17d5# => X"e0c42000",
		16#17d6# => X"e0631800",
		16#17d7# => X"9d66ffff",
		16#17d8# => X"e4862000",
		16#17d9# => X"10000003",
		16#17da# => X"9d000001",
		16#17db# => X"9d000000",
		16#17dc# => X"e0681800",
		16#17dd# => X"9ce00001",
		16#17de# => X"e48b3000",
		16#17df# => X"9d03ffff",
		16#17e0# => X"a8860000",
		16#17e1# => X"10000003",
		16#17e2# => X"9c42ffff",
		16#17e3# => X"9ce00000",
		16#17e4# => X"e0e74000",
		16#17e5# => X"19000fff",
		16#17e6# => X"a908ffff",
		16#17e7# => X"e4474000",
		16#17e8# => X"0fffffeb",
		16#17e9# => X"e4274000",
		16#17ea# => X"d405180c",
		16#17eb# => X"d4053010",
		16#17ec# => X"d4051008",
		16#17ed# => X"19a01fff",
		16#17ee# => X"9c400003",
		16#17ef# => X"a9adffff",
		16#17f0# => X"e4436800",
		16#17f1# => X"0c00000d",
		16#17f2# => X"d4051000",
		16#17f3# => X"b8e3001f",
		16#17f4# => X"b8440041",
		16#17f5# => X"84c50008",
		16#17f6# => X"a4840001",
		16#17f7# => X"e0471004",
		16#17f8# => X"b8630041",
		16#17f9# => X"e0441004",
		16#17fa# => X"9cc60001",
		16#17fb# => X"d405180c",
		16#17fc# => X"d4051010",
		16#17fd# => X"d4053008",
		16#17fe# => X"a9650000",
		16#17ff# => X"9c210008",
		16#1800# => X"8441fff8",
		16#1801# => X"44004800",
		16#1802# => X"85c1fffc",
		16#1803# => X"10000026",
		16#1804# => X"15000000",
		16#1805# => X"850b0004",
		16#1806# => X"84840004",
		16#1807# => X"9c400000",
		16#1808# => X"e4082000",
		16#1809# => X"0fffffa8",
		16#180a# => X"9c600000",
		16#180b# => X"e0833800",
		16#180c# => X"d4054004",
		16#180d# => X"d4056008",
		16#180e# => X"e4841800",
		16#180f# => X"10000003",
		16#1810# => X"9d000001",
		16#1811# => X"9d000000",
		16#1812# => X"e0423000",
		16#1813# => X"d4052010",
		16#1814# => X"e0681000",
		16#1815# => X"03ffffd8",
		16#1816# => X"d405180c",
		16#1817# => X"bc220002",
		16#1818# => X"13ffffe7",
		16#1819# => X"15000000",
		16#181a# => X"d4051000",
		16#181b# => X"844b0004",
		16#181c# => X"d4051004",
		16#181d# => X"844b0008",
		16#181e# => X"d4051008",
		16#181f# => X"844b000c",
		16#1820# => X"d405100c",
		16#1821# => X"844b0010",
		16#1822# => X"d4051010",
		16#1823# => X"844b0004",
		16#1824# => X"84640004",
		16#1825# => X"a9650000",
		16#1826# => X"e0431003",
		16#1827# => X"03ffffd8",
		16#1828# => X"d4051004",
		16#1829# => X"a98f0000",
		16#182a# => X"9cc00000",
		16#182b# => X"03ffff81",
		16#182c# => X"9ce00000",
		16#182d# => X"0fffffa8",
		16#182e# => X"15000000",
		16#182f# => X"03ffffbc",
		16#1830# => X"d405180c",
		16#1831# => X"e4443800",
		16#1832# => X"10000003",
		16#1833# => X"9d600001",
		16#1834# => X"a9680000",
		16#1835# => X"e0661002",
		16#1836# => X"e0635802",
		16#1837# => X"bd830000",
		16#1838# => X"0fffff87",
		16#1839# => X"9d600000",
		16#183a# => X"9c400001",
		16#183b# => X"e0802002",
		16#183c# => X"d4051004",
		16#183d# => X"bc440000",
		16#183e# => X"10000003",
		16#183f# => X"d4056008",
		16#1840# => X"9c400000",
		16#1841# => X"e0601802",
		16#1842# => X"d4052010",
		16#1843# => X"e0631002",
		16#1844# => X"03ffff7f",
		16#1845# => X"d405180c",
		16#1846# => X"9c210008",
		16#1847# => X"a9640000",
		16#1848# => X"8441fff8",
		16#1849# => X"44004800",
		16#184a# => X"85c1fffc",
		16#184b# => X"13ffff61",
		16#184c# => X"9da8ffe0",
		16#184d# => X"bd8d0000",
		16#184e# => X"1000002c",
		16#184f# => X"e18c4000",
		16#1850# => X"e1e66848",
		16#1851# => X"9ea00000",
		16#1852# => X"bd8d0000",
		16#1853# => X"10000024",
		16#1854# => X"9e200001",
		16#1855# => X"9d000000",
		16#1856# => X"e1b16808",
		16#1857# => X"9e28ffff",
		16#1858# => X"e4914000",
		16#1859# => X"10000003",
		16#185a# => X"9e600001",
		16#185b# => X"9e600000",
		16#185c# => X"9d0dffff",
		16#185d# => X"e2313803",
		16#185e# => X"e1134000",
		16#185f# => X"e1083003",
		16#1860# => X"a8d50000",
		16#1861# => X"e1088804",
		16#1862# => X"e1a04002",
		16#1863# => X"e10d4004",
		16#1864# => X"b908005f",
		16#1865# => X"03ffff47",
		16#1866# => X"e0e87804",
		16#1867# => X"9e20001f",
		16#1868# => X"ba6e0001",
		16#1869# => X"e2314002",
		16#186a# => X"e1e34048",
		16#186b# => X"e2338808",
		16#186c# => X"a9c20000",
		16#186d# => X"e1f17804",
		16#186e# => X"03ffff29",
		16#186f# => X"e2ae4048",
		16#1870# => X"0fffff61",
		16#1871# => X"15000000",
		16#1872# => X"03ffff7c",
		16#1873# => X"19a01fff",
		16#1874# => X"9da00000",
		16#1875# => X"03ffff27",
		16#1876# => X"e1114008",
		16#1877# => X"9da00000",
		16#1878# => X"03ffffdf",
		16#1879# => X"e1114008",
		16#187a# => X"9e20001f",
		16#187b# => X"ba660001",
		16#187c# => X"e2314002",
		16#187d# => X"e1e74048",
		16#187e# => X"e2338808",
		16#187f# => X"e2a64048",
		16#1880# => X"03ffffd2",
		16#1881# => X"e1f17804",
		16#1882# => X"bc230004",
		16#1883# => X"13ffff7c",
		16#1884# => X"15000000",
		16#1885# => X"846b0004",
		16#1886# => X"84440004",
		16#1887# => X"e4231000",
		16#1888# => X"0fffff77",
		16#1889# => X"15000000",
		16#188a# => X"19600001",
		16#188b# => X"03ffff74",
		16#188c# => X"a96b3d8c",
		16#188d# => X"d7e187ec",
		16#188e# => X"d7e14ffc",
		16#188f# => X"d7e117e4",
		16#1890# => X"d7e177e8",
		16#1891# => X"d7e197f0",
		16#1892# => X"d7e1a7f4",
		16#1893# => X"d7e1b7f8",
		16#1894# => X"84830000",
		16#1895# => X"9c21ffdc",
		16#1896# => X"8443000c",
		16#1897# => X"85c30010",
		16#1898# => X"bc440001",
		16#1899# => X"0c000051",
		16#189a# => X"86030004",
		16#189b# => X"bc040004",
		16#189c# => X"10000049",
		16#189d# => X"bc040002",
		16#189e# => X"1000002a",
		16#189f# => X"e0827004",
		16#18a0# => X"bc040000",
		16#18a1# => X"10000027",
		16#18a2# => X"15000000",
		16#18a3# => X"84630008",
		16#18a4# => X"bd63fc02",
		16#18a5# => X"0c00004e",
		16#18a6# => X"bd4303ff",
		16#18a7# => X"1000003e",
		16#18a8# => X"a48e00ff",
		16#18a9# => X"bc240080",
		16#18aa# => X"0c000031",
		16#18ab# => X"9c6303ff",
		16#18ac# => X"9c8e007f",
		16#18ad# => X"e4847000",
		16#18ae# => X"0c000035",
		16#18af# => X"9ca00001",
		16#18b0# => X"e0451000",
		16#18b1# => X"a9c40000",
		16#18b2# => X"18a01fff",
		16#18b3# => X"a8a5ffff",
		16#18b4# => X"e4422800",
		16#18b5# => X"0c000006",
		16#18b6# => X"b882001f",
		16#18b7# => X"b9ce0041",
		16#18b8# => X"b8420041",
		16#18b9# => X"9c630001",
		16#18ba# => X"e1c47004",
		16#18bb# => X"a4a307ff",
		16#18bc# => X"1900000f",
		16#18bd# => X"b8e20048",
		16#18be# => X"b8a50014",
		16#18bf# => X"a908ffff",
		16#18c0# => X"b8820018",
		16#18c1# => X"b9ce0048",
		16#18c2# => X"a8450000",
		16#18c3# => X"e0a74003",
		16#18c4# => X"9ce00000",
		16#18c5# => X"e0c47004",
		16#18c6# => X"00000006",
		16#18c7# => X"a8670000",
		16#18c8# => X"9c400000",
		16#18c9# => X"9c600000",
		16#18ca# => X"e0a20004",
		16#18cb# => X"e0c30004",
		16#18cc# => X"b890001f",
		16#18cd# => X"9c210024",
		16#18ce# => X"e0e51004",
		16#18cf# => X"8521fffc",
		16#18d0# => X"e0461804",
		16#18d1# => X"e0672004",
		16#18d2# => X"a9820000",
		16#18d3# => X"a9630000",
		16#18d4# => X"8441ffe4",
		16#18d5# => X"85c1ffe8",
		16#18d6# => X"8601ffec",
		16#18d7# => X"8641fff0",
		16#18d8# => X"8681fff4",
		16#18d9# => X"44004800",
		16#18da# => X"86c1fff8",
		16#18db# => X"a48e0100",
		16#18dc# => X"bc040000",
		16#18dd# => X"13ffffd6",
		16#18de# => X"18a01fff",
		16#18df# => X"9c8e0080",
		16#18e0# => X"e4847000",
		16#18e1# => X"13ffffcf",
		16#18e2# => X"9ca00001",
		16#18e3# => X"03ffffcd",
		16#18e4# => X"9ca00000",
		16#18e5# => X"18407ff0",
		16#18e6# => X"9c600000",
		16#18e7# => X"9ca00000",
		16#18e8# => X"03ffffe4",
		16#18e9# => X"9cc00000",
		16#18ea# => X"18600008",
		16#18eb# => X"1880000f",
		16#18ec# => X"e0421804",
		16#18ed# => X"a884ffff",
		16#18ee# => X"9c600000",
		16#18ef# => X"e0a22003",
		16#18f0# => X"a8ce0000",
		16#18f1# => X"03ffffdb",
		16#18f2# => X"18407ff0",
		16#18f3# => X"9e40fc02",
		16#18f4# => X"9ce00000",
		16#18f5# => X"9d000000",
		16#18f6# => X"e2521802",
		16#18f7# => X"d4013800",
		16#18f8# => X"d4014004",
		16#18f9# => X"bd520038",
		16#18fa# => X"10000046",
		16#18fb# => X"85010004",
		16#18fc# => X"a8620000",
		16#18fd# => X"a88e0000",
		16#18fe# => X"040004e6",
		16#18ff# => X"a8b20000",
		16#1900# => X"a8b20000",
		16#1901# => X"9c600000",
		16#1902# => X"9c800001",
		16#1903# => X"aacb0000",
		16#1904# => X"040004f4",
		16#1905# => X"aa8c0000",
		16#1906# => X"9c800001",
		16#1907# => X"a86b0000",
		16#1908# => X"bc2c0000",
		16#1909# => X"10000003",
		16#190a# => X"9cacffff",
		16#190b# => X"9c800000",
		16#190c# => X"9c63ffff",
		16#190d# => X"e1c57003",
		16#190e# => X"e0841800",
		16#190f# => X"d401b000",
		16#1910# => X"e0441003",
		16#1911# => X"e0427004",
		16#1912# => X"e0601002",
		16#1913# => X"e0431004",
		16#1914# => X"b842005f",
		16#1915# => X"e282a004",
		16#1916# => X"a45400ff",
		16#1917# => X"bc220080",
		16#1918# => X"10000027",
		16#1919# => X"d401a004",
		16#191a# => X"a4540100",
		16#191b# => X"bc020000",
		16#191c# => X"1000000e",
		16#191d# => X"85010000",
		16#191e# => X"9c540080",
		16#191f# => X"e482a000",
		16#1920# => X"0c000024",
		16#1921# => X"9c600001",
		16#1922# => X"84e10000",
		16#1923# => X"a8820000",
		16#1924# => X"e0a33800",
		16#1925# => X"a8640000",
		16#1926# => X"a8450000",
		16#1927# => X"d4011000",
		16#1928# => X"d4011804",
		16#1929# => X"85010000",
		16#192a# => X"84a10004",
		16#192b# => X"b8e80018",
		16#192c# => X"b8850048",
		16#192d# => X"b8480048",
		16#192e# => X"1900000f",
		16#192f# => X"e0c72004",
		16#1930# => X"18e00fff",
		16#1931# => X"a908ffff",
		16#1932# => X"84810000",
		16#1933# => X"a8e7ffff",
		16#1934# => X"e0a24003",
		16#1935# => X"e4443800",
		16#1936# => X"10000003",
		16#1937# => X"9c600001",
		16#1938# => X"9c600000",
		16#1939# => X"a48307ff",
		16#193a# => X"b8840014",
		16#193b# => X"a8440000",
		16#193c# => X"9c800000",
		16#193d# => X"03ffff8f",
		16#193e# => X"a8640000",
		16#193f# => X"85010004",
		16#1940# => X"9c48007f",
		16#1941# => X"e4824000",
		16#1942# => X"13ffffe0",
		16#1943# => X"9c600001",
		16#1944# => X"03ffffde",
		16#1945# => X"9c600000",
		16#1946# => X"d7e117fc",
		16#1947# => X"1840000f",
		16#1948# => X"84c30000",
		16#1949# => X"84a30004",
		16#194a# => X"b8e60054",
		16#194b# => X"b906005f",
		16#194c# => X"a842ffff",
		16#194d# => X"a4e707ff",
		16#194e# => X"d4044004",
		16#194f# => X"9c21fffc",
		16#1950# => X"bc270000",
		16#1951# => X"10000022",
		16#1952# => X"e0661003",
		16#1953# => X"e0c32804",
		16#1954# => X"bc260000",
		16#1955# => X"0c00002f",
		16#1956# => X"b8c50058",
		16#1957# => X"b8630008",
		16#1958# => X"9ce0fc02",
		16#1959# => X"b8a50008",
		16#195a# => X"e0661804",
		16#195b# => X"9cc00003",
		16#195c# => X"d4043808",
		16#195d# => X"d4043000",
		16#195e# => X"9cc0fc01",
		16#195f# => X"e0e52800",
		16#1960# => X"e0631800",
		16#1961# => X"e4872800",
		16#1962# => X"10000003",
		16#1963# => X"9d000001",
		16#1964# => X"9d000000",
		16#1965# => X"18400fff",
		16#1966# => X"e0681800",
		16#1967# => X"a842ffff",
		16#1968# => X"a9660000",
		16#1969# => X"a8a70000",
		16#196a# => X"e4431000",
		16#196b# => X"0ffffff4",
		16#196c# => X"9cc6ffff",
		16#196d# => X"9c210004",
		16#196e# => X"d4045808",
		16#196f# => X"d404180c",
		16#1970# => X"d4043810",
		16#1971# => X"44004800",
		16#1972# => X"8441fffc",
		16#1973# => X"bc2707ff",
		16#1974# => X"0c000015",
		16#1975# => X"9ce7fc01",
		16#1976# => X"b8c50058",
		16#1977# => X"b8630008",
		16#1978# => X"18401000",
		16#1979# => X"e0661804",
		16#197a# => X"b8a50008",
		16#197b# => X"e0631004",
		16#197c# => X"d4043808",
		16#197d# => X"9cc00003",
		16#197e# => X"d4043000",
		16#197f# => X"d404180c",
		16#1980# => X"d4042810",
		16#1981# => X"9c210004",
		16#1982# => X"44004800",
		16#1983# => X"8441fffc",
		16#1984# => X"9c600002",
		16#1985# => X"9c210004",
		16#1986# => X"d4041800",
		16#1987# => X"44004800",
		16#1988# => X"8441fffc",
		16#1989# => X"e0e32804",
		16#198a# => X"bc270000",
		16#198b# => X"0c00000a",
		16#198c# => X"15000000",
		16#198d# => X"18400008",
		16#198e# => X"e0c61003",
		16#198f# => X"bc060000",
		16#1990# => X"13ffffee",
		16#1991# => X"15000000",
		16#1992# => X"9cc00001",
		16#1993# => X"03ffffec",
		16#1994# => X"d4043000",
		16#1995# => X"9c600004",
		16#1996# => X"03ffffeb",
		16#1997# => X"d4041800",
		16#1998# => X"d7e14ffc",
		16#1999# => X"d7e117f4",
		16#199a# => X"d7e177f8",
		16#199b# => X"9c21ffa8",
		16#199c# => X"9dc10028",
		16#199d# => X"d4011844",
		16#199e# => X"d4012048",
		16#199f# => X"9c610044",
		16#19a0# => X"a88e0000",
		16#19a1# => X"d401283c",
		16#19a2# => X"d4013040",
		16#19a3# => X"07ffffa3",
		16#19a4# => X"9c410014",
		16#19a5# => X"9c61003c",
		16#19a6# => X"07ffffa0",
		16#19a7# => X"a8820000",
		16#19a8# => X"a86e0000",
		16#19a9# => X"a8820000",
		16#19aa# => X"07fffdc4",
		16#19ab# => X"a8a10000",
		16#19ac# => X"07fffee1",
		16#19ad# => X"a86b0000",
		16#19ae# => X"9c210058",
		16#19af# => X"a84b0000",
		16#19b0# => X"a86c0000",
		16#19b1# => X"8521fffc",
		16#19b2# => X"e1620004",
		16#19b3# => X"e1830004",
		16#19b4# => X"85c1fff8",
		16#19b5# => X"44004800",
		16#19b6# => X"8441fff4",
		16#19b7# => X"d7e14ffc",
		16#19b8# => X"d7e117f4",
		16#19b9# => X"d7e177f8",
		16#19ba# => X"9c21ffa8",
		16#19bb# => X"9c410028",
		16#19bc# => X"d4011844",
		16#19bd# => X"d4012048",
		16#19be# => X"9c610044",
		16#19bf# => X"a8820000",
		16#19c0# => X"d401283c",
		16#19c1# => X"d4013040",
		16#19c2# => X"07ffff84",
		16#19c3# => X"9dc10014",
		16#19c4# => X"9c61003c",
		16#19c5# => X"07ffff81",
		16#19c6# => X"a88e0000",
		16#19c7# => X"84c10018",
		16#19c8# => X"a88e0000",
		16#19c9# => X"acc60001",
		16#19ca# => X"a8a10000",
		16#19cb# => X"a8620000",
		16#19cc# => X"07fffda2",
		16#19cd# => X"d4013018",
		16#19ce# => X"07fffebf",
		16#19cf# => X"a86b0000",
		16#19d0# => X"9c210058",
		16#19d1# => X"a84b0000",
		16#19d2# => X"a86c0000",
		16#19d3# => X"8521fffc",
		16#19d4# => X"e1620004",
		16#19d5# => X"e1830004",
		16#19d6# => X"85c1fff8",
		16#19d7# => X"44004800",
		16#19d8# => X"8441fff4",
		16#19d9# => X"d7e14ffc",
		16#19da# => X"d7e117dc",
		16#19db# => X"d7e177e0",
		16#19dc# => X"d7e187e4",
		16#19dd# => X"d7e197e8",
		16#19de# => X"d7e1a7ec",
		16#19df# => X"d7e1b7f0",
		16#19e0# => X"d7e1c7f4",
		16#19e1# => X"d7e1d7f8",
		16#19e2# => X"9c21ff90",
		16#19e3# => X"9dc10028",
		16#19e4# => X"d4011844",
		16#19e5# => X"d4012048",
		16#19e6# => X"9c610044",
		16#19e7# => X"a88e0000",
		16#19e8# => X"d401283c",
		16#19e9# => X"d4013040",
		16#19ea# => X"07ffff5c",
		16#19eb# => X"9e010014",
		16#19ec# => X"9c61003c",
		16#19ed# => X"07ffff59",
		16#19ee# => X"a8900000",
		16#19ef# => X"84410028",
		16#19f0# => X"bc420001",
		16#19f1# => X"0c0000c7",
		16#19f2# => X"84a10014",
		16#19f3# => X"bc450001",
		16#19f4# => X"0c0000df",
		16#19f5# => X"bc220004",
		16#19f6# => X"0c0000be",
		16#19f7# => X"bc250004",
		16#19f8# => X"0c0000d7",
		16#19f9# => X"bc220002",
		16#19fa# => X"0c0000be",
		16#19fb# => X"bc250002",
		16#19fc# => X"0c0000d7",
		16#19fd# => X"84410038",
		16#19fe# => X"9c600000",
		16#19ff# => X"86010024",
		16#1a00# => X"a8a30000",
		16#1a01# => X"a8820000",
		16#1a02# => X"a8d00000",
		16#1a03# => X"040003c4",
		16#1a04# => X"86810020",
		16#1a05# => X"9c600000",
		16#1a06# => X"a8940000",
		16#1a07# => X"a8a30000",
		16#1a08# => X"a8c20000",
		16#1a09# => X"a9cb0000",
		16#1a0a# => X"040003bd",
		16#1a0b# => X"ab0c0000",
		16#1a0c# => X"9c600000",
		16#1a0d# => X"87410034",
		16#1a0e# => X"a8a30000",
		16#1a0f# => X"a8d40000",
		16#1a10# => X"a89a0000",
		16#1a11# => X"aa4c0000",
		16#1a12# => X"040003b5",
		16#1a13# => X"a84b0000",
		16#1a14# => X"9c600000",
		16#1a15# => X"a89a0000",
		16#1a16# => X"a8a30000",
		16#1a17# => X"a8d00000",
		16#1a18# => X"aa8b0000",
		16#1a19# => X"040003ae",
		16#1a1a# => X"aacc0000",
		16#1a1b# => X"e0ac9000",
		16#1a1c# => X"a90b0000",
		16#1a1d# => X"e4856000",
		16#1a1e# => X"0c00006d",
		16#1a1f# => X"9da00001",
		16#1a20# => X"e0e81000",
		16#1a21# => X"e0ed3800",
		16#1a22# => X"e4423800",
		16#1a23# => X"0c000063",
		16#1a24# => X"e4223800",
		16#1a25# => X"9c400001",
		16#1a26# => X"9c600000",
		16#1a27# => X"e0a57000",
		16#1a28# => X"e44e2800",
		16#1a29# => X"0c000009",
		16#1a2a# => X"a8d80000",
		16#1a2b# => X"9c830001",
		16#1a2c# => X"e4841800",
		16#1a2d# => X"0c000081",
		16#1a2e# => X"9d000001",
		16#1a2f# => X"e1081000",
		16#1a30# => X"a8640000",
		16#1a31# => X"a8480000",
		16#1a32# => X"e187b000",
		16#1a33# => X"e48c3800",
		16#1a34# => X"10000003",
		16#1a35# => X"9c800001",
		16#1a36# => X"9c800000",
		16#1a37# => X"e10c1800",
		16#1a38# => X"e084a000",
		16#1a39# => X"e4886000",
		16#1a3a# => X"10000003",
		16#1a3b# => X"9da00001",
		16#1a3c# => X"9da00000",
		16#1a3d# => X"84e10018",
		16#1a3e# => X"8581002c",
		16#1a3f# => X"85c1001c",
		16#1a40# => X"e18c3805",
		16#1a41# => X"84e10030",
		16#1a42# => X"e1606002",
		16#1a43# => X"e0ee3800",
		16#1a44# => X"e18b6004",
		16#1a45# => X"e0841000",
		16#1a46# => X"b98c005f",
		16#1a47# => X"9c670004",
		16#1a48# => X"18401fff",
		16#1a49# => X"e08d2000",
		16#1a4a# => X"d4011808",
		16#1a4b# => X"a842ffff",
		16#1a4c# => X"d4016004",
		16#1a4d# => X"e4441000",
		16#1a4e# => X"0c000017",
		16#1a4f# => X"a8680000",
		16#1a50# => X"9ce70005",
		16#1a51# => X"b9030041",
		16#1a52# => X"a4630001",
		16#1a53# => X"b964001f",
		16#1a54# => X"b985001f",
		16#1a55# => X"b8460041",
		16#1a56# => X"b9a50041",
		16#1a57# => X"b8840041",
		16#1a58# => X"bc030000",
		16#1a59# => X"10000005",
		16#1a5a# => X"a9e70000",
		16#1a5b# => X"18608000",
		16#1a5c# => X"e0cc1004",
		16#1a5d# => X"e0ad1804",
		16#1a5e# => X"e06b4004",
		16#1a5f# => X"19001fff",
		16#1a60# => X"a908ffff",
		16#1a61# => X"e4444000",
		16#1a62# => X"13ffffef",
		16#1a63# => X"9ce70001",
		16#1a64# => X"d4017808",
		16#1a65# => X"19600fff",
		16#1a66# => X"a96bffff",
		16#1a67# => X"e4445800",
		16#1a68# => X"1000002c",
		16#1a69# => X"84e10008",
		16#1a6a# => X"0000000d",
		16#1a6b# => X"e1631800",
		16#1a6c# => X"e4883000",
		16#1a6d# => X"10000003",
		16#1a6e# => X"9ca00001",
		16#1a6f# => X"9ca00000",
		16#1a70# => X"18400fff",
		16#1a71# => X"a8c80000",
		16#1a72# => X"a842ffff",
		16#1a73# => X"e44b1000",
		16#1a74# => X"1000001f",
		16#1a75# => X"e0a56800",
		16#1a76# => X"e1631800",
		16#1a77# => X"e0842000",
		16#1a78# => X"e1063000",
		16#1a79# => X"e1a52800",
		16#1a7a# => X"9d800001",
		16#1a7b# => X"e48b1800",
		16#1a7c# => X"10000003",
		16#1a7d# => X"9ce7ffff",
		16#1a7e# => X"9d800000",
		16#1a7f# => X"e08c2000",
		16#1a80# => X"a86b0000",
		16#1a81# => X"bd850000",
		16#1a82# => X"0fffffea",
		16#1a83# => X"a9640000",
		16#1a84# => X"03ffffe8",
		16#1a85# => X"a8630001",
		16#1a86# => X"0c00002a",
		16#1a87# => X"e4522800",
		16#1a88# => X"9c400000",
		16#1a89# => X"03ffff9e",
		16#1a8a# => X"9c600000",
		16#1a8b# => X"9da00000",
		16#1a8c# => X"e0e81000",
		16#1a8d# => X"e0ed3800",
		16#1a8e# => X"e4423800",
		16#1a8f# => X"13ffff96",
		16#1a90# => X"e4223800",
		16#1a91# => X"03fffff5",
		16#1a92# => X"15000000",
		16#1a93# => X"d4013808",
		16#1a94# => X"a44300ff",
		16#1a95# => X"bc220080",
		16#1a96# => X"0c00002b",
		16#1a97# => X"a4430100",
		16#1a98# => X"9c400003",
		16#1a99# => X"d4011810",
		16#1a9a# => X"d401200c",
		16#1a9b# => X"d4011000",
		16#1a9c# => X"a8610000",
		16#1a9d# => X"07fffdf0",
		16#1a9e# => X"15000000",
		16#1a9f# => X"9c210070",
		16#1aa0# => X"a84b0000",
		16#1aa1# => X"a86c0000",
		16#1aa2# => X"8521fffc",
		16#1aa3# => X"e1620004",
		16#1aa4# => X"e1830004",
		16#1aa5# => X"85c1ffe0",
		16#1aa6# => X"8441ffdc",
		16#1aa7# => X"8601ffe4",
		16#1aa8# => X"8641ffe8",
		16#1aa9# => X"8681ffec",
		16#1aaa# => X"86c1fff0",
		16#1aab# => X"8701fff4",
		16#1aac# => X"44004800",
		16#1aad# => X"8741fff8",
		16#1aae# => X"03ffff81",
		16#1aaf# => X"9d000000",
		16#1ab0# => X"13ffff75",
		16#1ab1# => X"9c400000",
		16#1ab2# => X"03ffff75",
		16#1ab3# => X"9c600000",
		16#1ab4# => X"18600001",
		16#1ab5# => X"bc050002",
		16#1ab6# => X"13ffffe7",
		16#1ab7# => X"a8633d8c",
		16#1ab8# => X"8481002c",
		16#1ab9# => X"84410018",
		16#1aba# => X"a86e0000",
		16#1abb# => X"e0441005",
		16#1abc# => X"e0801002",
		16#1abd# => X"e0441004",
		16#1abe# => X"b842005f",
		16#1abf# => X"03ffffde",
		16#1ac0# => X"d401102c",
		16#1ac1# => X"bc220000",
		16#1ac2# => X"13ffffd6",
		16#1ac3# => X"e0a53004",
		16#1ac4# => X"bc050000",
		16#1ac5# => X"13ffffd3",
		16#1ac6# => X"9ca30080",
		16#1ac7# => X"e4851800",
		16#1ac8# => X"10000003",
		16#1ac9# => X"9cc00001",
		16#1aca# => X"a8c20000",
		16#1acb# => X"9ce0ff00",
		16#1acc# => X"e0862000",
		16#1acd# => X"03ffffcb",
		16#1ace# => X"e0653803",
		16#1acf# => X"18600001",
		16#1ad0# => X"bc020002",
		16#1ad1# => X"13ffffcc",
		16#1ad2# => X"a8633d8c",
		16#1ad3# => X"84410018",
		16#1ad4# => X"8481002c",
		16#1ad5# => X"a8700000",
		16#1ad6# => X"e0441005",
		16#1ad7# => X"e0801002",
		16#1ad8# => X"e0441004",
		16#1ad9# => X"b842005f",
		16#1ada# => X"03ffffc3",
		16#1adb# => X"d4011018",
		16#1adc# => X"d7e14ffc",
		16#1add# => X"d7e117f0",
		16#1ade# => X"d7e177f4",
		16#1adf# => X"d7e187f8",
		16#1ae0# => X"9c21ffb8",
		16#1ae1# => X"9dc10014",
		16#1ae2# => X"d4011830",
		16#1ae3# => X"d4012034",
		16#1ae4# => X"9c610030",
		16#1ae5# => X"d4012828",
		16#1ae6# => X"d401302c",
		16#1ae7# => X"07fffe5f",
		16#1ae8# => X"a88e0000",
		16#1ae9# => X"9c610028",
		16#1aea# => X"07fffe5c",
		16#1aeb# => X"a8810000",
		16#1aec# => X"84410014",
		16#1aed# => X"bca20001",
		16#1aee# => X"10000059",
		16#1aef# => X"a86e0000",
		16#1af0# => X"84a10000",
		16#1af1# => X"bca50001",
		16#1af2# => X"10000055",
		16#1af3# => X"a8610000",
		16#1af4# => X"84810018",
		16#1af5# => X"84610004",
		16#1af6# => X"bc020004",
		16#1af7# => X"e0641805",
		16#1af8# => X"10000063",
		16#1af9# => X"d4011818",
		16#1afa# => X"bc220002",
		16#1afb# => X"0c000060",
		16#1afc# => X"bc250004",
		16#1afd# => X"0c000080",
		16#1afe# => X"bc250002",
		16#1aff# => X"0c00007a",
		16#1b00# => X"84410008",
		16#1b01# => X"8461001c",
		16#1b02# => X"84c10020",
		16#1b03# => X"e0431002",
		16#1b04# => X"8621000c",
		16#1b05# => X"d401101c",
		16#1b06# => X"84a10024",
		16#1b07# => X"e4513000",
		16#1b08# => X"0c00004b",
		16#1b09# => X"86e10010",
		16#1b0a# => X"e0652800",
		16#1b0b# => X"e4832800",
		16#1b0c# => X"0c000055",
		16#1b0d# => X"9c800001",
		16#1b0e# => X"e0c63000",
		16#1b0f# => X"9c42ffff",
		16#1b10# => X"e0c43000",
		16#1b11# => X"a8a30000",
		16#1b12# => X"d401101c",
		16#1b13# => X"9da0003d",
		16#1b14# => X"18401000",
		16#1b15# => X"9c600000",
		16#1b16# => X"9d600000",
		16#1b17# => X"9d800000",
		16#1b18# => X"baa2001f",
		16#1b19# => X"b9e30041",
		16#1b1a# => X"ba620041",
		16#1b1b# => X"9dadffff",
		16#1b1c# => X"e1f57804",
		16#1b1d# => X"a8f30000",
		16#1b1e# => X"e4513000",
		16#1b1f# => X"10000015",
		16#1b20# => X"a90f0000",
		16#1b21# => X"e1eb1004",
		16#1b22# => X"e2ac1804",
		16#1b23# => X"a84f0000",
		16#1b24# => X"e2668802",
		16#1b25# => X"e1e5b802",
		16#1b26# => X"e4313000",
		16#1b27# => X"10000005",
		16#1b28# => X"a8750000",
		16#1b29# => X"e4572800",
		16#1b2a# => X"1000000a",
		16#1b2b# => X"15000000",
		16#1b2c# => X"e44f2800",
		16#1b2d# => X"9cc00001",
		16#1b2e# => X"e1620004",
		16#1b2f# => X"e1830004",
		16#1b30# => X"10000003",
		16#1b31# => X"a8af0000",
		16#1b32# => X"9cc00000",
		16#1b33# => X"e0d33002",
		16#1b34# => X"e1e52800",
		16#1b35# => X"e0c63000",
		16#1b36# => X"e48f2800",
		16#1b37# => X"e0470004",
		16#1b38# => X"e0680004",
		16#1b39# => X"10000003",
		16#1b3a# => X"9e600001",
		16#1b3b# => X"9e600000",
		16#1b3c# => X"a8af0000",
		16#1b3d# => X"bc2d0000",
		16#1b3e# => X"13ffffda",
		16#1b3f# => X"e0d33000",
		16#1b40# => X"a46c00ff",
		16#1b41# => X"bc230080",
		16#1b42# => X"0c000026",
		16#1b43# => X"a88b0000",
		16#1b44# => X"a86e0000",
		16#1b45# => X"d4015820",
		16#1b46# => X"d4016024",
		16#1b47# => X"07fffd46",
		16#1b48# => X"15000000",
		16#1b49# => X"9c210048",
		16#1b4a# => X"a84b0000",
		16#1b4b# => X"a86c0000",
		16#1b4c# => X"8521fffc",
		16#1b4d# => X"e1620004",
		16#1b4e# => X"e1830004",
		16#1b4f# => X"85c1fff4",
		16#1b50# => X"8441fff0",
		16#1b51# => X"44004800",
		16#1b52# => X"8601fff8",
		16#1b53# => X"e4313000",
		16#1b54# => X"13ffffc0",
		16#1b55# => X"9da0003d",
		16#1b56# => X"e4572800",
		16#1b57# => X"0fffffbd",
		16#1b58# => X"e0652800",
		16#1b59# => X"03ffffb3",
		16#1b5a# => X"e4832800",
		16#1b5b# => X"18600001",
		16#1b5c# => X"e4022800",
		16#1b5d# => X"13ffffea",
		16#1b5e# => X"a8633d8c",
		16#1b5f# => X"03ffffe8",
		16#1b60# => X"a86e0000",
		16#1b61# => X"9c800000",
		16#1b62# => X"e0c63000",
		16#1b63# => X"9c42ffff",
		16#1b64# => X"e0c43000",
		16#1b65# => X"a8a30000",
		16#1b66# => X"03ffffad",
		16#1b67# => X"d401101c",
		16#1b68# => X"a46c0100",
		16#1b69# => X"bc230000",
		16#1b6a# => X"13ffffdb",
		16#1b6b# => X"a86e0000",
		16#1b6c# => X"e0c67804",
		16#1b6d# => X"bc060000",
		16#1b6e# => X"13ffffd7",
		16#1b6f# => X"15000000",
		16#1b70# => X"9c6c0080",
		16#1b71# => X"e4836000",
		16#1b72# => X"10000003",
		16#1b73# => X"9ca00001",
		16#1b74# => X"a8ad0000",
		16#1b75# => X"9c40ff00",
		16#1b76# => X"e1652000",
		16#1b77# => X"03ffffcd",
		16#1b78# => X"e1831003",
		16#1b79# => X"9c400004",
		16#1b7a# => X"a86e0000",
		16#1b7b# => X"03ffffcc",
		16#1b7c# => X"d4011014",
		16#1b7d# => X"9c600000",
		16#1b7e# => X"9c400000",
		16#1b7f# => X"d4011020",
		16#1b80# => X"d4011824",
		16#1b81# => X"9c600000",
		16#1b82# => X"d401181c",
		16#1b83# => X"03ffffc4",
		16#1b84# => X"a86e0000",
		16#1b85# => X"84a30000",
		16#1b86# => X"9d600001",
		16#1b87# => X"e4a55800",
		16#1b88# => X"10000016",
		16#1b89# => X"15000000",
		16#1b8a# => X"84c40000",
		16#1b8b# => X"e4a65800",
		16#1b8c# => X"10000012",
		16#1b8d# => X"bc250004",
		16#1b8e# => X"0c000044",
		16#1b8f# => X"bc260004",
		16#1b90# => X"0c000019",
		16#1b91# => X"bc250002",
		16#1b92# => X"0c000014",
		16#1b93# => X"bc260002",
		16#1b94# => X"0c00000c",
		16#1b95# => X"15000000",
		16#1b96# => X"84a30004",
		16#1b97# => X"84c40004",
		16#1b98# => X"e4053000",
		16#1b99# => X"10000016",
		16#1b9a# => X"15000000",
		16#1b9b# => X"bc050000",
		16#1b9c# => X"0c000008",
		16#1b9d# => X"15000000",
		16#1b9e# => X"44004800",
		16#1b9f# => X"15000000",
		16#1ba0# => X"84630004",
		16#1ba1# => X"bc030000",
		16#1ba2# => X"13fffffc",
		16#1ba3# => X"15000000",
		16#1ba4# => X"44004800",
		16#1ba5# => X"9d60ffff",
		16#1ba6# => X"bc060002",
		16#1ba7# => X"13fffff7",
		16#1ba8# => X"9d600000",
		16#1ba9# => X"84640004",
		16#1baa# => X"bc030000",
		16#1bab# => X"13fffff3",
		16#1bac# => X"9d60ffff",
		16#1bad# => X"44004800",
		16#1bae# => X"9d600001",
		16#1baf# => X"84e30008",
		16#1bb0# => X"84c40008",
		16#1bb1# => X"e5a73000",
		16#1bb2# => X"0fffffea",
		16#1bb3# => X"bc050000",
		16#1bb4# => X"e5673000",
		16#1bb5# => X"0c000015",
		16#1bb6# => X"bc050000",
		16#1bb7# => X"84c3000c",
		16#1bb8# => X"84e4000c",
		16#1bb9# => X"84630010",
		16#1bba# => X"e4463800",
		16#1bbb# => X"10000013",
		16#1bbc# => X"84840010",
		16#1bbd# => X"e4263800",
		16#1bbe# => X"10000005",
		16#1bbf# => X"e4473000",
		16#1bc0# => X"e4432000",
		16#1bc1# => X"1000000d",
		16#1bc2# => X"e4473000",
		16#1bc3# => X"10000007",
		16#1bc4# => X"bc050000",
		16#1bc5# => X"e4273000",
		16#1bc6# => X"1000000a",
		16#1bc7# => X"e4441800",
		16#1bc8# => X"0c000008",
		16#1bc9# => X"bc050000",
		16#1bca# => X"0fffffe3",
		16#1bcb# => X"9d60ffff",
		16#1bcc# => X"44004800",
		16#1bcd# => X"15000000",
		16#1bce# => X"03ffffcd",
		16#1bcf# => X"9d600001",
		16#1bd0# => X"44004800",
		16#1bd1# => X"9d600000",
		16#1bd2# => X"13ffffce",
		16#1bd3# => X"15000000",
		16#1bd4# => X"85640004",
		16#1bd5# => X"84630004",
		16#1bd6# => X"44004800",
		16#1bd7# => X"e16b1802",
		16#1bd8# => X"d7e14ffc",
		16#1bd9# => X"d7e117f4",
		16#1bda# => X"d7e177f8",
		16#1bdb# => X"9c21ffbc",
		16#1bdc# => X"9dc10014",
		16#1bdd# => X"d4011830",
		16#1bde# => X"d4012034",
		16#1bdf# => X"9c610030",
		16#1be0# => X"d4012828",
		16#1be1# => X"d401302c",
		16#1be2# => X"07fffd64",
		16#1be3# => X"a88e0000",
		16#1be4# => X"9c610028",
		16#1be5# => X"07fffd61",
		16#1be6# => X"a8810000",
		16#1be7# => X"a86e0000",
		16#1be8# => X"07ffff9d",
		16#1be9# => X"a8810000",
		16#1bea# => X"9c210044",
		16#1beb# => X"8521fffc",
		16#1bec# => X"8441fff4",
		16#1bed# => X"44004800",
		16#1bee# => X"85c1fff8",
		16#1bef# => X"d7e14ffc",
		16#1bf0# => X"d7e177f8",
		16#1bf1# => X"d7e117f4",
		16#1bf2# => X"9c21ffbc",
		16#1bf3# => X"9dc10014",
		16#1bf4# => X"d4011830",
		16#1bf5# => X"d4012034",
		16#1bf6# => X"9c610030",
		16#1bf7# => X"d4012828",
		16#1bf8# => X"d401302c",
		16#1bf9# => X"07fffd4d",
		16#1bfa# => X"a88e0000",
		16#1bfb# => X"9c610028",
		16#1bfc# => X"07fffd4a",
		16#1bfd# => X"a8810000",
		16#1bfe# => X"9d600001",
		16#1bff# => X"84610014",
		16#1c00# => X"e4a35800",
		16#1c01# => X"10000007",
		16#1c02# => X"84610000",
		16#1c03# => X"e4a35800",
		16#1c04# => X"10000004",
		16#1c05# => X"a86e0000",
		16#1c06# => X"07ffff7f",
		16#1c07# => X"a8810000",
		16#1c08# => X"9c210044",
		16#1c09# => X"8521fffc",
		16#1c0a# => X"8441fff4",
		16#1c0b# => X"44004800",
		16#1c0c# => X"85c1fff8",
		16#1c0d# => X"d7e14ffc",
		16#1c0e# => X"d7e177f8",
		16#1c0f# => X"d7e117f4",
		16#1c10# => X"9c21ffbc",
		16#1c11# => X"9dc10014",
		16#1c12# => X"d4011830",
		16#1c13# => X"d4012034",
		16#1c14# => X"9c610030",
		16#1c15# => X"d4012828",
		16#1c16# => X"d401302c",
		16#1c17# => X"07fffd2f",
		16#1c18# => X"a88e0000",
		16#1c19# => X"9c610028",
		16#1c1a# => X"07fffd2c",
		16#1c1b# => X"a8810000",
		16#1c1c# => X"9d600001",
		16#1c1d# => X"84610014",
		16#1c1e# => X"e4a35800",
		16#1c1f# => X"10000007",
		16#1c20# => X"84610000",
		16#1c21# => X"e4a35800",
		16#1c22# => X"10000004",
		16#1c23# => X"a86e0000",
		16#1c24# => X"07ffff61",
		16#1c25# => X"a8810000",
		16#1c26# => X"9c210044",
		16#1c27# => X"8521fffc",
		16#1c28# => X"8441fff4",
		16#1c29# => X"44004800",
		16#1c2a# => X"85c1fff8",
		16#1c2b# => X"d7e14ffc",
		16#1c2c# => X"d7e177f8",
		16#1c2d# => X"d7e117f4",
		16#1c2e# => X"9c21ffbc",
		16#1c2f# => X"9dc10014",
		16#1c30# => X"d4011830",
		16#1c31# => X"d4012034",
		16#1c32# => X"9c610030",
		16#1c33# => X"d4012828",
		16#1c34# => X"d401302c",
		16#1c35# => X"07fffd11",
		16#1c36# => X"a88e0000",
		16#1c37# => X"9c610028",
		16#1c38# => X"07fffd0e",
		16#1c39# => X"a8810000",
		16#1c3a# => X"84610014",
		16#1c3b# => X"bca30001",
		16#1c3c# => X"10000008",
		16#1c3d# => X"9d60ffff",
		16#1c3e# => X"84610000",
		16#1c3f# => X"bca30001",
		16#1c40# => X"10000004",
		16#1c41# => X"a86e0000",
		16#1c42# => X"07ffff43",
		16#1c43# => X"a8810000",
		16#1c44# => X"9c210044",
		16#1c45# => X"8521fffc",
		16#1c46# => X"8441fff4",
		16#1c47# => X"44004800",
		16#1c48# => X"85c1fff8",
		16#1c49# => X"d7e14ffc",
		16#1c4a# => X"d7e177f8",
		16#1c4b# => X"d7e117f4",
		16#1c4c# => X"9c21ffbc",
		16#1c4d# => X"9dc10014",
		16#1c4e# => X"d4011830",
		16#1c4f# => X"d4012034",
		16#1c50# => X"9c610030",
		16#1c51# => X"d4012828",
		16#1c52# => X"d401302c",
		16#1c53# => X"07fffcf3",
		16#1c54# => X"a88e0000",
		16#1c55# => X"9c610028",
		16#1c56# => X"07fffcf0",
		16#1c57# => X"a8810000",
		16#1c58# => X"84610014",
		16#1c59# => X"bca30001",
		16#1c5a# => X"10000008",
		16#1c5b# => X"9d60ffff",
		16#1c5c# => X"84610000",
		16#1c5d# => X"bca30001",
		16#1c5e# => X"10000004",
		16#1c5f# => X"a86e0000",
		16#1c60# => X"07ffff25",
		16#1c61# => X"a8810000",
		16#1c62# => X"9c210044",
		16#1c63# => X"8521fffc",
		16#1c64# => X"8441fff4",
		16#1c65# => X"44004800",
		16#1c66# => X"85c1fff8",
		16#1c67# => X"d7e14ffc",
		16#1c68# => X"d7e177f8",
		16#1c69# => X"d7e117f4",
		16#1c6a# => X"9c21ffbc",
		16#1c6b# => X"9dc10014",
		16#1c6c# => X"d4011830",
		16#1c6d# => X"d4012034",
		16#1c6e# => X"9c610030",
		16#1c6f# => X"d4012828",
		16#1c70# => X"d401302c",
		16#1c71# => X"07fffcd5",
		16#1c72# => X"a88e0000",
		16#1c73# => X"9c610028",
		16#1c74# => X"07fffcd2",
		16#1c75# => X"a8810000",
		16#1c76# => X"9d600001",
		16#1c77# => X"84610014",
		16#1c78# => X"e4a35800",
		16#1c79# => X"10000007",
		16#1c7a# => X"84610000",
		16#1c7b# => X"e4a35800",
		16#1c7c# => X"10000004",
		16#1c7d# => X"a86e0000",
		16#1c7e# => X"07ffff07",
		16#1c7f# => X"a8810000",
		16#1c80# => X"9c210044",
		16#1c81# => X"8521fffc",
		16#1c82# => X"8441fff4",
		16#1c83# => X"44004800",
		16#1c84# => X"85c1fff8",
		16#1c85# => X"d7e14ffc",
		16#1c86# => X"d7e177f8",
		16#1c87# => X"d7e117f4",
		16#1c88# => X"9c21ffbc",
		16#1c89# => X"9dc10014",
		16#1c8a# => X"d4011830",
		16#1c8b# => X"d4012034",
		16#1c8c# => X"9c610030",
		16#1c8d# => X"d4012828",
		16#1c8e# => X"d401302c",
		16#1c8f# => X"07fffcb7",
		16#1c90# => X"a88e0000",
		16#1c91# => X"9c610028",
		16#1c92# => X"07fffcb4",
		16#1c93# => X"a8810000",
		16#1c94# => X"9d600001",
		16#1c95# => X"84610014",
		16#1c96# => X"e4a35800",
		16#1c97# => X"10000007",
		16#1c98# => X"84610000",
		16#1c99# => X"e4a35800",
		16#1c9a# => X"10000004",
		16#1c9b# => X"a86e0000",
		16#1c9c# => X"07fffee9",
		16#1c9d# => X"a8810000",
		16#1c9e# => X"9c210044",
		16#1c9f# => X"8521fffc",
		16#1ca0# => X"8441fff4",
		16#1ca1# => X"44004800",
		16#1ca2# => X"85c1fff8",
		16#1ca3# => X"d7e14ffc",
		16#1ca4# => X"9c21ffc4",
		16#1ca5# => X"d4011830",
		16#1ca6# => X"d4012034",
		16#1ca7# => X"9c610030",
		16#1ca8# => X"d4012828",
		16#1ca9# => X"d401302c",
		16#1caa# => X"07fffc9c",
		16#1cab# => X"9c810014",
		16#1cac# => X"9c610028",
		16#1cad# => X"07fffc99",
		16#1cae# => X"a8810000",
		16#1caf# => X"9d600001",
		16#1cb0# => X"84610014",
		16#1cb1# => X"e4a35800",
		16#1cb2# => X"10000005",
		16#1cb3# => X"84610000",
		16#1cb4# => X"e4a35800",
		16#1cb5# => X"0c000006",
		16#1cb6# => X"15000000",
		16#1cb7# => X"9c21003c",
		16#1cb8# => X"8521fffc",
		16#1cb9# => X"44004800",
		16#1cba# => X"15000000",
		16#1cbb# => X"9c21003c",
		16#1cbc# => X"8521fffc",
		16#1cbd# => X"44004800",
		16#1cbe# => X"9d600000",
		16#1cbf# => X"b883005f",
		16#1cc0# => X"d7e117f8",
		16#1cc1# => X"d7e14ffc",
		16#1cc2# => X"9c400003",
		16#1cc3# => X"9c21ffe4",
		16#1cc4# => X"bc230000",
		16#1cc5# => X"d4011000",
		16#1cc6# => X"1000000a",
		16#1cc7# => X"d4012004",
		16#1cc8# => X"9c400002",
		16#1cc9# => X"d4011000",
		16#1cca# => X"07fffbc3",
		16#1ccb# => X"a8610000",
		16#1ccc# => X"9c21001c",
		16#1ccd# => X"8521fffc",
		16#1cce# => X"44004800",
		16#1ccf# => X"8441fff8",
		16#1cd0# => X"a8430000",
		16#1cd1# => X"9c60003c",
		16#1cd2# => X"bc040000",
		16#1cd3# => X"0c000015",
		16#1cd4# => X"d4011808",
		16#1cd5# => X"9c800000",
		16#1cd6# => X"a8620000",
		16#1cd7# => X"d401200c",
		16#1cd8# => X"04000134",
		16#1cd9# => X"d4011010",
		16#1cda# => X"9c8b001d",
		16#1cdb# => X"bda40000",
		16#1cdc# => X"13ffffee",
		16#1cdd# => X"9d6bfffd",
		16#1cde# => X"bd8b0000",
		16#1cdf# => X"1000000f",
		16#1ce0# => X"e1625808",
		16#1ce1# => X"9c400000",
		16#1ce2# => X"d401580c",
		16#1ce3# => X"d4011010",
		16#1ce4# => X"9c40003c",
		16#1ce5# => X"e0822002",
		16#1ce6# => X"03ffffe4",
		16#1ce7# => X"d4012008",
		16#1ce8# => X"18608000",
		16#1ce9# => X"e4021800",
		16#1cea# => X"1000000c",
		16#1ceb# => X"1960c1e0",
		16#1cec# => X"03ffffe9",
		16#1ced# => X"e0401002",
		16#1cee# => X"9ca0001f",
		16#1cef# => X"b8620041",
		16#1cf0# => X"e0a52002",
		16#1cf1# => X"e0422008",
		16#1cf2# => X"e0a32848",
		16#1cf3# => X"d4011010",
		16#1cf4# => X"03fffff0",
		16#1cf5# => X"d401280c",
		16#1cf6# => X"03ffffd6",
		16#1cf7# => X"9d800000",
		16#1cf8# => X"d7e117f8",
		16#1cf9# => X"9c800000",
		16#1cfa# => X"d7e14ffc",
		16#1cfb# => X"9c21ffe4",
		16#1cfc# => X"a8430000",
		16#1cfd# => X"e4232000",
		16#1cfe# => X"0c000023",
		16#1cff# => X"d4012004",
		16#1d00# => X"9c800003",
		16#1d01# => X"9ca00000",
		16#1d02# => X"d4012000",
		16#1d03# => X"9c80003c",
		16#1d04# => X"d4011810",
		16#1d05# => X"d4012008",
		16#1d06# => X"04000106",
		16#1d07# => X"d401280c",
		16#1d08# => X"9c6b001d",
		16#1d09# => X"bd630000",
		16#1d0a# => X"0c00001a",
		16#1d0b# => X"bc030000",
		16#1d0c# => X"1000000b",
		16#1d0d# => X"9d6bfffd",
		16#1d0e# => X"bd8b0000",
		16#1d0f# => X"1000002a",
		16#1d10# => X"e1625808",
		16#1d11# => X"9c400000",
		16#1d12# => X"d401580c",
		16#1d13# => X"d4011010",
		16#1d14# => X"9c40003c",
		16#1d15# => X"e0621802",
		16#1d16# => X"d4011808",
		16#1d17# => X"07fffb76",
		16#1d18# => X"a8610000",
		16#1d19# => X"9c21001c",
		16#1d1a# => X"a84b0000",
		16#1d1b# => X"a86c0000",
		16#1d1c# => X"8521fffc",
		16#1d1d# => X"e1620004",
		16#1d1e# => X"e1830004",
		16#1d1f# => X"44004800",
		16#1d20# => X"8441fff8",
		16#1d21# => X"9c400002",
		16#1d22# => X"03fffff5",
		16#1d23# => X"d4011000",
		16#1d24# => X"e0801802",
		16#1d25# => X"9cc4ffe0",
		16#1d26# => X"bd860000",
		16#1d27# => X"1000001a",
		16#1d28# => X"9ca00000",
		16#1d29# => X"9ca5ffff",
		16#1d2a# => X"e0822048",
		16#1d2b# => X"e0a51003",
		16#1d2c# => X"b8c6009f",
		16#1d2d# => X"e0402802",
		16#1d2e# => X"e0a22804",
		16#1d2f# => X"e0843003",
		16#1d30# => X"b845005f",
		16#1d31# => X"9ca0003c",
		16#1d32# => X"e0422004",
		16#1d33# => X"e0651802",
		16#1d34# => X"9ca00000",
		16#1d35# => X"d4011808",
		16#1d36# => X"d401280c",
		16#1d37# => X"03ffffe0",
		16#1d38# => X"d4011010",
		16#1d39# => X"9c80001f",
		16#1d3a# => X"b8a20041",
		16#1d3b# => X"e0841802",
		16#1d3c# => X"e0421808",
		16#1d3d# => X"e0852048",
		16#1d3e# => X"d4011010",
		16#1d3f# => X"03ffffd5",
		16#1d40# => X"d401200c",
		16#1d41# => X"9ca00001",
		16#1d42# => X"03ffffe7",
		16#1d43# => X"e0a52008",
		16#1d44# => X"d7e14ffc",
		16#1d45# => X"9c21ffe0",
		16#1d46# => X"d4011814",
		16#1d47# => X"d4012018",
		16#1d48# => X"9c610014",
		16#1d49# => X"07fffbfd",
		16#1d4a# => X"a8810000",
		16#1d4b# => X"84610000",
		16#1d4c# => X"bc030002",
		16#1d4d# => X"10000018",
		16#1d4e# => X"9d600000",
		16#1d4f# => X"bca30001",
		16#1d50# => X"10000015",
		16#1d51# => X"bc230004",
		16#1d52# => X"0c000020",
		16#1d53# => X"84610008",
		16#1d54# => X"bd830000",
		16#1d55# => X"10000010",
		16#1d56# => X"bda3001e",
		16#1d57# => X"0c000012",
		16#1d58# => X"9d60003c",
		16#1d59# => X"e06b1802",
		16#1d5a# => X"9c83ffe0",
		16#1d5b# => X"bd840000",
		16#1d5c# => X"1000001e",
		16#1d5d# => X"84a1000c",
		16#1d5e# => X"8561000c",
		16#1d5f# => X"e16b2048",
		16#1d60# => X"84610004",
		16#1d61# => X"bc030000",
		16#1d62# => X"10000003",
		16#1d63# => X"15000000",
		16#1d64# => X"e1605802",
		16#1d65# => X"9c210020",
		16#1d66# => X"8521fffc",
		16#1d67# => X"44004800",
		16#1d68# => X"15000000",
		16#1d69# => X"84610004",
		16#1d6a# => X"bc030000",
		16#1d6b# => X"0c00000b",
		16#1d6c# => X"15000000",
		16#1d6d# => X"9c210020",
		16#1d6e# => X"19607fff",
		16#1d6f# => X"8521fffc",
		16#1d70# => X"44004800",
		16#1d71# => X"a96bffff",
		16#1d72# => X"84610004",
		16#1d73# => X"e4035800",
		16#1d74# => X"13fffff9",
		16#1d75# => X"15000000",
		16#1d76# => X"9c210020",
		16#1d77# => X"8521fffc",
		16#1d78# => X"44004800",
		16#1d79# => X"19608000",
		16#1d7a# => X"9c80001f",
		16#1d7b# => X"b8a50001",
		16#1d7c# => X"e0841802",
		16#1d7d# => X"85610010",
		16#1d7e# => X"e0852008",
		16#1d7f# => X"e16b1848",
		16#1d80# => X"03ffffe0",
		16#1d81# => X"e1645804",
		16#1d82# => X"d7e14ffc",
		16#1d83# => X"d7e117f8",
		16#1d84# => X"9c21ffdc",
		16#1d85# => X"d4011814",
		16#1d86# => X"d4012018",
		16#1d87# => X"9c610014",
		16#1d88# => X"07fffbbe",
		16#1d89# => X"a8810000",
		16#1d8a# => X"84810004",
		16#1d8b# => X"a8610000",
		16#1d8c# => X"e0402002",
		16#1d8d# => X"e0422004",
		16#1d8e# => X"ac42ffff",
		16#1d8f# => X"b842005f",
		16#1d90# => X"07fffafd",
		16#1d91# => X"d4011004",
		16#1d92# => X"9c210024",
		16#1d93# => X"a84b0000",
		16#1d94# => X"a86c0000",
		16#1d95# => X"8521fffc",
		16#1d96# => X"e1620004",
		16#1d97# => X"e1830004",
		16#1d98# => X"44004800",
		16#1d99# => X"8441fff8",
		16#1d9a# => X"d7e14ffc",
		16#1d9b# => X"d7e117f8",
		16#1d9c# => X"9c21ffe4",
		16#1d9d# => X"d4011800",
		16#1d9e# => X"d4012004",
		16#1d9f# => X"d4012808",
		16#1da0# => X"d401300c",
		16#1da1# => X"d4013810",
		16#1da2# => X"07fffaeb",
		16#1da3# => X"a8610000",
		16#1da4# => X"9c21001c",
		16#1da5# => X"a84b0000",
		16#1da6# => X"a86c0000",
		16#1da7# => X"8521fffc",
		16#1da8# => X"e1620004",
		16#1da9# => X"e1830004",
		16#1daa# => X"44004800",
		16#1dab# => X"8441fff8",
		16#1dac# => X"d7e117f8",
		16#1dad# => X"d7e14ffc",
		16#1dae# => X"9c21ffdc",
		16#1daf# => X"18403fff",
		16#1db0# => X"d4011814",
		16#1db1# => X"d4012018",
		16#1db2# => X"9c610014",
		16#1db3# => X"a8810000",
		16#1db4# => X"07fffb92",
		16#1db5# => X"a842ffff",
		16#1db6# => X"84610010",
		16#1db7# => X"84c1000c",
		16#1db8# => X"b883005e",
		16#1db9# => X"b8c60002",
		16#1dba# => X"e0631003",
		16#1dbb# => X"bc030000",
		16#1dbc# => X"10000003",
		16#1dbd# => X"e0c62004",
		16#1dbe# => X"a8c60001",
		16#1dbf# => X"84610000",
		16#1dc0# => X"84810004",
		16#1dc1# => X"07fff98b",
		16#1dc2# => X"84a10008",
		16#1dc3# => X"9c210024",
		16#1dc4# => X"8521fffc",
		16#1dc5# => X"44004800",
		16#1dc6# => X"8441fff8",
		16#1dc7# => X"a4e4ffff",
		16#1dc8# => X"b9040050",
		16#1dc9# => X"a566ffff",
		16#1dca# => X"b9860050",
		16#1dcb# => X"e1ab3b06",
		16#1dcc# => X"e16b4306",
		16#1dcd# => X"e0ec3b06",
		16#1dce# => X"b9ed0050",
		16#1dcf# => X"e0eb3800",
		16#1dd0# => X"d7e117fc",
		16#1dd1# => X"e0e77800",
		16#1dd2# => X"9c21fffc",
		16#1dd3# => X"e4ab3800",
		16#1dd4# => X"10000004",
		16#1dd5# => X"e10c4306",
		16#1dd6# => X"18400001",
		16#1dd7# => X"e1081000",
		16#1dd8# => X"e0c61b06",
		16#1dd9# => X"e0842b06",
		16#1dda# => X"b8670050",
		16#1ddb# => X"b8e70010",
		16#1ddc# => X"a5adffff",
		16#1ddd# => X"e1081800",
		16#1dde# => X"e1643000",
		16#1ddf# => X"9c210004",
		16#1de0# => X"e1876800",
		16#1de1# => X"e16b4000",
		16#1de2# => X"44004800",
		16#1de3# => X"8441fffc",
		16#1de4# => X"bc050000",
		16#1de5# => X"1000000b",
		16#1de6# => X"9cc00020",
		16#1de7# => X"e0c62802",
		16#1de8# => X"bd460000",
		16#1de9# => X"0c00000a",
		16#1dea# => X"15000000",
		16#1deb# => X"e0c33008",
		16#1dec# => X"e0842848",
		16#1ded# => X"e0a32848",
		16#1dee# => X"e0862004",
		16#1def# => X"a8650000",
		16#1df0# => X"a9630000",
		16#1df1# => X"44004800",
		16#1df2# => X"a9840000",
		16#1df3# => X"e0803002",
		16#1df4# => X"9ca00000",
		16#1df5# => X"e0832048",
		16#1df6# => X"03fffffa",
		16#1df7# => X"a8650000",
		16#1df8# => X"bc050000",
		16#1df9# => X"1000000b",
		16#1dfa# => X"9cc00020",
		16#1dfb# => X"e0c62802",
		16#1dfc# => X"bd460000",
		16#1dfd# => X"0c00000a",
		16#1dfe# => X"15000000",
		16#1dff# => X"e0c43048",
		16#1e00# => X"e0632808",
		16#1e01# => X"e0a42808",
		16#1e02# => X"e0661804",
		16#1e03# => X"a8850000",
		16#1e04# => X"a9630000",
		16#1e05# => X"44004800",
		16#1e06# => X"a9840000",
		16#1e07# => X"e0603002",
		16#1e08# => X"9ca00000",
		16#1e09# => X"e0641808",
		16#1e0a# => X"03fffffa",
		16#1e0b# => X"a8850000",
		16#1e0c# => X"d7e117fc",
		16#1e0d# => X"a840ffff",
		16#1e0e# => X"e4431000",
		16#1e0f# => X"10000010",
		16#1e10# => X"9c21fffc",
		16#1e11# => X"bc4300ff",
		16#1e12# => X"0c000018",
		16#1e13# => X"9c800020",
		16#1e14# => X"9c800018",
		16#1e15# => X"9ca00008",
		16#1e16# => X"18400001",
		16#1e17# => X"e0632848",
		16#1e18# => X"a8423da0",
		16#1e19# => X"9c210004",
		16#1e1a# => X"e0631000",
		16#1e1b# => X"8441fffc",
		16#1e1c# => X"8d630000",
		16#1e1d# => X"44004800",
		16#1e1e# => X"e1645802",
		16#1e1f# => X"184000ff",
		16#1e20# => X"a842ffff",
		16#1e21# => X"e4431000",
		16#1e22# => X"10000005",
		16#1e23# => X"15000000",
		16#1e24# => X"9c800010",
		16#1e25# => X"03fffff1",
		16#1e26# => X"a8a40000",
		16#1e27# => X"9c800008",
		16#1e28# => X"03ffffee",
		16#1e29# => X"9ca00018",
		16#1e2a# => X"03ffffec",
		16#1e2b# => X"9ca00000",
		16#1e2c# => X"d7e14ffc",
		16#1e2d# => X"9c21fffc",
		16#1e2e# => X"a8830000",
		16#1e2f# => X"9c210004",
		16#1e30# => X"9c600000",
		16#1e31# => X"8521fffc",
		16#1e32# => X"a8a30000",
		16#1e33# => X"00001018",
		16#1e34# => X"a8c30000",
		16#1e35# => X"d7e117f8",
		16#1e36# => X"d7e14ffc",
		16#1e37# => X"9c800000",
		16#1e38# => X"9c21fff8",
		16#1e39# => X"04001063",
		16#1e3a# => X"a8430000",
		16#1e3b# => X"18800001",
		16#1e3c# => X"a8843ea0",
		16#1e3d# => X"84840000",
		16#1e3e# => X"84a4003c",
		16#1e3f# => X"bc050000",
		16#1e40# => X"10000004",
		16#1e41# => X"15000000",
		16#1e42# => X"48002800",
		16#1e43# => X"a8640000",
		16#1e44# => X"04002e4d",
		16#1e45# => X"a8620000",
		16#1e46# => X"a8830000",
		16#1e47# => X"18600001",
		16#1e48# => X"d7e14ffc",
		16#1e49# => X"a86363e0",
		16#1e4a# => X"9c21fffc",
		16#1e4b# => X"84630000",
		16#1e4c# => X"9c210004",
		16#1e4d# => X"8521fffc",
		16#1e4e# => X"0000000c",
		16#1e4f# => X"15000000",
		16#1e50# => X"a8830000",
		16#1e51# => X"18600001",
		16#1e52# => X"d7e14ffc",
		16#1e53# => X"a86363e0",
		16#1e54# => X"9c21fffc",
		16#1e55# => X"84630000",
		16#1e56# => X"9c210004",
		16#1e57# => X"8521fffc",
		16#1e58# => X"00001ab7",
		16#1e59# => X"15000000",
		16#1e5a# => X"d7e177dc",
		16#1e5b# => X"d7e187e0",
		16#1e5c# => X"d7e14ffc",
		16#1e5d# => X"d7e117d8",
		16#1e5e# => X"d7e197e4",
		16#1e5f# => X"d7e1a7e8",
		16#1e60# => X"d7e1b7ec",
		16#1e61# => X"d7e1c7f0",
		16#1e62# => X"d7e1d7f4",
		16#1e63# => X"d7e1e7f8",
		16#1e64# => X"9dc4000b",
		16#1e65# => X"9c21ffd8",
		16#1e66# => X"bcae0016",
		16#1e67# => X"10000036",
		16#1e68# => X"aa030000",
		16#1e69# => X"9c40fff8",
		16#1e6a# => X"e1ce1003",
		16#1e6b# => X"b86e005f",
		16#1e6c# => X"e48e2000",
		16#1e6d# => X"10000003",
		16#1e6e# => X"9c400001",
		16#1e6f# => X"9c400000",
		16#1e70# => X"a44200ff",
		16#1e71# => X"bc220000",
		16#1e72# => X"100000b3",
		16#1e73# => X"bc030000",
		16#1e74# => X"0c0000b2",
		16#1e75# => X"9c40000c",
		16#1e76# => X"04000234",
		16#1e77# => X"a8700000",
		16#1e78# => X"bc4e01f7",
		16#1e79# => X"10000027",
		16#1e7a# => X"b8ee0049",
		16#1e7b# => X"18800001",
		16#1e7c# => X"b8ee0043",
		16#1e7d# => X"a8846808",
		16#1e7e# => X"e06e2000",
		16#1e7f# => X"8443000c",
		16#1e80# => X"e4221800",
		16#1e81# => X"0c00018e",
		16#1e82# => X"aa440000",
		16#1e83# => X"84820004",
		16#1e84# => X"9ca0fffc",
		16#1e85# => X"8462000c",
		16#1e86# => X"e0842803",
		16#1e87# => X"84c20008",
		16#1e88# => X"e0822000",
		16#1e89# => X"d406180c",
		16#1e8a# => X"84a40004",
		16#1e8b# => X"d4033008",
		16#1e8c# => X"a8a50001",
		16#1e8d# => X"a8700000",
		16#1e8e# => X"0400021e",
		16#1e8f# => X"d4042804",
		16#1e90# => X"9d620008",
		16#1e91# => X"9c210028",
		16#1e92# => X"8521fffc",
		16#1e93# => X"8441ffd8",
		16#1e94# => X"85c1ffdc",
		16#1e95# => X"8601ffe0",
		16#1e96# => X"8641ffe4",
		16#1e97# => X"8681ffe8",
		16#1e98# => X"86c1ffec",
		16#1e99# => X"8701fff0",
		16#1e9a# => X"8741fff4",
		16#1e9b# => X"44004800",
		16#1e9c# => X"8781fff8",
		16#1e9d# => X"9c600000",
		16#1e9e# => X"03ffffce",
		16#1e9f# => X"9dc00010",
		16#1ea0# => X"bc270000",
		16#1ea1# => X"0c000088",
		16#1ea2# => X"bc470004",
		16#1ea3# => X"10000155",
		16#1ea4# => X"bc470014",
		16#1ea5# => X"b8ee0046",
		16#1ea6# => X"9ce70038",
		16#1ea7# => X"b8670003",
		16#1ea8# => X"19600001",
		16#1ea9# => X"a96b6808",
		16#1eaa# => X"e0635800",
		16#1eab# => X"8443000c",
		16#1eac# => X"e4031000",
		16#1ead# => X"10000019",
		16#1eae# => X"aa4b0000",
		16#1eaf# => X"9ca0fffc",
		16#1eb0# => X"84820004",
		16#1eb1# => X"e0842803",
		16#1eb2# => X"e0a47002",
		16#1eb3# => X"bd45000f",
		16#1eb4# => X"100000b9",
		16#1eb5# => X"bd650000",
		16#1eb6# => X"0c00000c",
		16#1eb7# => X"15000000",
		16#1eb8# => X"000000b8",
		16#1eb9# => X"e0822000",
		16#1eba# => X"84820004",
		16#1ebb# => X"e0845803",
		16#1ebc# => X"e0a47002",
		16#1ebd# => X"bda5000f",
		16#1ebe# => X"0c0000af",
		16#1ebf# => X"bd850000",
		16#1ec0# => X"0c0000af",
		16#1ec1# => X"15000000",
		16#1ec2# => X"8442000c",
		16#1ec3# => X"e4231000",
		16#1ec4# => X"13fffff6",
		16#1ec5# => X"9d60fffc",
		16#1ec6# => X"9ce70001",
		16#1ec7# => X"18c00001",
		16#1ec8# => X"a8c66810",
		16#1ec9# => X"84460008",
		16#1eca# => X"e4261000",
		16#1ecb# => X"0c00007f",
		16#1ecc# => X"9c60fffc",
		16#1ecd# => X"84820004",
		16#1ece# => X"e0841803",
		16#1ecf# => X"e0647002",
		16#1ed0# => X"bda3000f",
		16#1ed1# => X"0c00012f",
		16#1ed2# => X"bd830000",
		16#1ed3# => X"d406300c",
		16#1ed4# => X"0c0000a7",
		16#1ed5# => X"d4063008",
		16#1ed6# => X"bc4401ff",
		16#1ed7# => X"10000055",
		16#1ed8# => X"b8640049",
		16#1ed9# => X"b8640043",
		16#1eda# => X"9d000001",
		16#1edb# => X"84920004",
		16#1edc# => X"b8a30082",
		16#1edd# => X"b8630003",
		16#1ede# => X"e1082808",
		16#1edf# => X"18a00001",
		16#1ee0# => X"a8a56808",
		16#1ee1# => X"e0882004",
		16#1ee2# => X"e0632800",
		16#1ee3# => X"d4122004",
		16#1ee4# => X"84a30008",
		16#1ee5# => X"d402180c",
		16#1ee6# => X"d4022808",
		16#1ee7# => X"d4031008",
		16#1ee8# => X"d405100c",
		16#1ee9# => X"b8470082",
		16#1eea# => X"9c600001",
		16#1eeb# => X"e0631008",
		16#1eec# => X"e4432000",
		16#1eed# => X"10000064",
		16#1eee# => X"e0441803",
		16#1eef# => X"bc220000",
		16#1ef0# => X"1000000d",
		16#1ef1# => X"9c40fffc",
		16#1ef2# => X"e0631800",
		16#1ef3# => X"e0e71003",
		16#1ef4# => X"e0441803",
		16#1ef5# => X"bc220000",
		16#1ef6# => X"10000007",
		16#1ef7# => X"9ce70004",
		16#1ef8# => X"e0631800",
		16#1ef9# => X"e0432003",
		16#1efa# => X"bc020000",
		16#1efb# => X"13fffffd",
		16#1efc# => X"9ce70004",
		16#1efd# => X"18800001",
		16#1efe# => X"b9870003",
		16#1eff# => X"a8846808",
		16#1f00# => X"a9670000",
		16#1f01# => X"e18c2000",
		16#1f02# => X"a90c0000",
		16#1f03# => X"8448000c",
		16#1f04# => X"e4081000",
		16#1f05# => X"10000019",
		16#1f06# => X"9c80fffc",
		16#1f07# => X"84a20004",
		16#1f08# => X"e0a52003",
		16#1f09# => X"e0857002",
		16#1f0a# => X"bd44000f",
		16#1f0b# => X"1000010b",
		16#1f0c# => X"bd640000",
		16#1f0d# => X"0c00000d",
		16#1f0e# => X"15000000",
		16#1f0f# => X"0000011b",
		16#1f10# => X"e0a22800",
		16#1f11# => X"9c80fffc",
		16#1f12# => X"84a20004",
		16#1f13# => X"e0a52003",
		16#1f14# => X"e0857002",
		16#1f15# => X"bda4000f",
		16#1f16# => X"0c000100",
		16#1f17# => X"bd840000",
		16#1f18# => X"0c000111",
		16#1f19# => X"15000000",
		16#1f1a# => X"8442000c",
		16#1f1b# => X"e4281000",
		16#1f1c# => X"13fffff5",
		16#1f1d# => X"15000000",
		16#1f1e# => X"9d6b0001",
		16#1f1f# => X"a44b0003",
		16#1f20# => X"bc220000",
		16#1f21# => X"0c000142",
		16#1f22# => X"9d080008",
		16#1f23# => X"03ffffe1",
		16#1f24# => X"8448000c",
		16#1f25# => X"9c40000c",
		16#1f26# => X"9d600000",
		16#1f27# => X"03ffff6a",
		16#1f28# => X"d4101000",
		16#1f29# => X"b8ee0043",
		16#1f2a# => X"03ffff7e",
		16#1f2b# => X"b8670003",
		16#1f2c# => X"bc430004",
		16#1f2d# => X"1000010b",
		16#1f2e# => X"bc430014",
		16#1f2f# => X"b9040046",
		16#1f30# => X"9d080038",
		16#1f31# => X"19600001",
		16#1f32# => X"b8a80003",
		16#1f33# => X"a96b6808",
		16#1f34# => X"e0a55800",
		16#1f35# => X"84650008",
		16#1f36# => X"e4032800",
		16#1f37# => X"0c000008",
		16#1f38# => X"b9080082",
		16#1f39# => X"00000114",
		16#1f3a# => X"9c800001",
		16#1f3b# => X"84630008",
		16#1f3c# => X"e4051800",
		16#1f3d# => X"10000008",
		16#1f3e# => X"15000000",
		16#1f3f# => X"85030004",
		16#1f40# => X"9d60fffc",
		16#1f41# => X"e1085803",
		16#1f42# => X"e4844000",
		16#1f43# => X"13fffff8",
		16#1f44# => X"15000000",
		16#1f45# => X"8483000c",
		16#1f46# => X"d402200c",
		16#1f47# => X"d4021808",
		16#1f48# => X"d4041008",
		16#1f49# => X"d403100c",
		16#1f4a# => X"b8470082",
		16#1f4b# => X"9c600001",
		16#1f4c# => X"84920004",
		16#1f4d# => X"e0631008",
		16#1f4e# => X"e4432000",
		16#1f4f# => X"0fffffa0",
		16#1f50# => X"e0441803",
		16#1f51# => X"84520008",
		16#1f52# => X"9ca0fffc",
		16#1f53# => X"86820004",
		16#1f54# => X"e2942803",
		16#1f55# => X"e0747002",
		16#1f56# => X"bda3000f",
		16#1f57# => X"10000003",
		16#1f58# => X"9c800001",
		16#1f59# => X"9c800000",
		16#1f5a# => X"a48400ff",
		16#1f5b# => X"bc240000",
		16#1f5c# => X"10000027",
		16#1f5d# => X"e44ea000",
		16#1f5e# => X"0c0000de",
		16#1f5f# => X"9ca00001",
		16#1f60# => X"a4a500ff",
		16#1f61# => X"bc050000",
		16#1f62# => X"0c000021",
		16#1f63# => X"a88e0001",
		16#1f64# => X"a8630001",
		16#1f65# => X"e1c27000",
		16#1f66# => X"d4022004",
		16#1f67# => X"d40e1804",
		16#1f68# => X"d4127008",
		16#1f69# => X"04000143",
		16#1f6a# => X"a8700000",
		16#1f6b# => X"03ffff26",
		16#1f6c# => X"9d620008",
		16#1f6d# => X"03ffff59",
		16#1f6e# => X"9ce7ffff",
		16#1f6f# => X"e0822000",
		16#1f70# => X"8462000c",
		16#1f71# => X"84a40004",
		16#1f72# => X"84c20008",
		16#1f73# => X"a8a50001",
		16#1f74# => X"d406180c",
		16#1f75# => X"d4033008",
		16#1f76# => X"d4042804",
		16#1f77# => X"04000135",
		16#1f78# => X"a8700000",
		16#1f79# => X"03ffff18",
		16#1f7a# => X"9d620008",
		16#1f7b# => X"e0822000",
		16#1f7c# => X"a8700000",
		16#1f7d# => X"84a40004",
		16#1f7e# => X"a8a50001",
		16#1f7f# => X"0400012d",
		16#1f80# => X"d4042804",
		16#1f81# => X"03ffff10",
		16#1f82# => X"9d620008",
		16#1f83# => X"18600001",
		16#1f84# => X"1b800001",
		16#1f85# => X"a8637a78",
		16#1f86# => X"ab9c6c14",
		16#1f87# => X"86c30000",
		16#1f88# => X"847c0000",
		16#1f89# => X"9ed60010",
		16#1f8a# => X"bc03ffff",
		16#1f8b# => X"10000005",
		16#1f8c# => X"e2d67000",
		16#1f8d# => X"9ed60fff",
		16#1f8e# => X"9d60f000",
		16#1f8f# => X"e2d65803",
		16#1f90# => X"a8700000",
		16#1f91# => X"040005af",
		16#1f92# => X"a8960000",
		16#1f93# => X"bc2bffff",
		16#1f94# => X"0c0000ec",
		16#1f95# => X"ab0b0000",
		16#1f96# => X"e082a000",
		16#1f97# => X"e4a45800",
		16#1f98# => X"0c0000a6",
		16#1f99# => X"18a00001",
		16#1f9a# => X"1b400001",
		16#1f9b# => X"e4245800",
		16#1f9c# => X"ab5a7a84",
		16#1f9d# => X"847a0000",
		16#1f9e# => X"e0761800",
		16#1f9f# => X"0c0000eb",
		16#1fa0# => X"d41a1800",
		16#1fa1# => X"84bc0000",
		16#1fa2# => X"bc25ffff",
		16#1fa3# => X"0c0000f9",
		16#1fa4# => X"e06b1800",
		16#1fa5# => X"e0832002",
		16#1fa6# => X"d41a2000",
		16#1fa7# => X"a46b0007",
		16#1fa8# => X"bc030000",
		16#1fa9# => X"10000006",
		16#1faa# => X"9c801000",
		16#1fab# => X"9c800008",
		16#1fac# => X"e0641802",
		16#1fad# => X"e30b1800",
		16#1fae# => X"9c831000",
		16#1faf# => X"e2d8b000",
		16#1fb0# => X"a8700000",
		16#1fb1# => X"a6d60fff",
		16#1fb2# => X"e2c4b002",
		16#1fb3# => X"0400058d",
		16#1fb4# => X"a8960000",
		16#1fb5# => X"bc0bffff",
		16#1fb6# => X"100000e4",
		16#1fb7# => X"9c800001",
		16#1fb8# => X"e08bc002",
		16#1fb9# => X"e084b000",
		16#1fba# => X"a8840001",
		16#1fbb# => X"847a0000",
		16#1fbc# => X"d4182004",
		16#1fbd# => X"e0761800",
		16#1fbe# => X"18800001",
		16#1fbf# => X"d412c008",
		16#1fc0# => X"a8846808",
		16#1fc1# => X"e4022000",
		16#1fc2# => X"10000011",
		16#1fc3# => X"d41a1800",
		16#1fc4# => X"bc54000f",
		16#1fc5# => X"0c000099",
		16#1fc6# => X"9ca0fff8",
		16#1fc7# => X"9c94fff4",
		16#1fc8# => X"9cc00005",
		16#1fc9# => X"e0842803",
		16#1fca# => X"e0a22000",
		16#1fcb# => X"bca4000f",
		16#1fcc# => X"d4053004",
		16#1fcd# => X"d4053008",
		16#1fce# => X"84a20004",
		16#1fcf# => X"a4a50001",
		16#1fd0# => X"e0842804",
		16#1fd1# => X"0c0000c2",
		16#1fd2# => X"d4022004",
		16#1fd3# => X"18400001",
		16#1fd4# => X"a8427a7c",
		16#1fd5# => X"84820000",
		16#1fd6# => X"e4a32000",
		16#1fd7# => X"10000003",
		16#1fd8# => X"18800001",
		16#1fd9# => X"d4021800",
		16#1fda# => X"a8847a80",
		16#1fdb# => X"84440000",
		16#1fdc# => X"e4431000",
		16#1fdd# => X"0c000065",
		16#1fde# => X"15000000",
		16#1fdf# => X"d4041800",
		16#1fe0# => X"84520008",
		16#1fe1# => X"9c60fffc",
		16#1fe2# => X"84820004",
		16#1fe3# => X"e0841803",
		16#1fe4# => X"e0647002",
		16#1fe5# => X"bda3000f",
		16#1fe6# => X"10000003",
		16#1fe7# => X"9ca00001",
		16#1fe8# => X"9ca00000",
		16#1fe9# => X"a4a500ff",
		16#1fea# => X"bc250000",
		16#1feb# => X"10000009",
		16#1fec# => X"e44e2000",
		16#1fed# => X"10000003",
		16#1fee# => X"9cc00001",
		16#1fef# => X"a8c50000",
		16#1ff0# => X"a4c600ff",
		16#1ff1# => X"bc060000",
		16#1ff2# => X"13ffff72",
		16#1ff3# => X"a88e0001",
		16#1ff4# => X"040000b8",
		16#1ff5# => X"a8700000",
		16#1ff6# => X"03fffe9b",
		16#1ff7# => X"9d600000",
		16#1ff8# => X"0c00003d",
		16#1ff9# => X"bc470054",
		16#1ffa# => X"1000004d",
		16#1ffb# => X"bc470154",
		16#1ffc# => X"b8ee004c",
		16#1ffd# => X"9ce7006e",
		16#1ffe# => X"03fffeaa",
		16#1fff# => X"b8670003",
		16#2000# => X"e0827000",
		16#2001# => X"a9ce0001",
		16#2002# => X"a8e30001",
		16#2003# => X"e0a41800",
		16#2004# => X"d4027004",
		16#2005# => X"d406200c",
		16#2006# => X"d4062008",
		16#2007# => X"d4051800",
		16#2008# => X"d404300c",
		16#2009# => X"d4043008",
		16#200a# => X"d4043804",
		16#200b# => X"040000a1",
		16#200c# => X"a8700000",
		16#200d# => X"03fffe84",
		16#200e# => X"9d620008",
		16#200f# => X"9c620008",
		16#2010# => X"8443000c",
		16#2011# => X"e4031000",
		16#2012# => X"0ffffe71",
		16#2013# => X"9ce70002",
		16#2014# => X"03fffeb4",
		16#2015# => X"18c00001",
		16#2016# => X"e0627000",
		16#2017# => X"84a2000c",
		16#2018# => X"84e20008",
		16#2019# => X"a9ce0001",
		16#201a# => X"d407280c",
		16#201b# => X"d4053808",
		16#201c# => X"e0a32000",
		16#201d# => X"a8e40001",
		16#201e# => X"d406180c",
		16#201f# => X"d4061808",
		16#2020# => X"d4027004",
		16#2021# => X"d403300c",
		16#2022# => X"d4033008",
		16#2023# => X"d4033804",
		16#2024# => X"d4052000",
		16#2025# => X"04000087",
		16#2026# => X"a8700000",
		16#2027# => X"03fffe6a",
		16#2028# => X"9d620008",
		16#2029# => X"e0a22800",
		16#202a# => X"8462000c",
		16#202b# => X"84c50004",
		16#202c# => X"84820008",
		16#202d# => X"a8c60001",
		16#202e# => X"d404180c",
		16#202f# => X"d4032008",
		16#2030# => X"d4053004",
		16#2031# => X"0400007b",
		16#2032# => X"a8700000",
		16#2033# => X"03fffe5e",
		16#2034# => X"9d620008",
		16#2035# => X"9ce7005b",
		16#2036# => X"03fffe72",
		16#2037# => X"b8670003",
		16#2038# => X"10000021",
		16#2039# => X"bc430054",
		16#203a# => X"03fffef7",
		16#203b# => X"9d03005b",
		16#203c# => X"03ffff24",
		16#203d# => X"a8a40000",
		16#203e# => X"a8a56808",
		16#203f# => X"e4022800",
		16#2040# => X"13ffff5a",
		16#2041# => X"15000000",
		16#2042# => X"84520008",
		16#2043# => X"9d60fffc",
		16#2044# => X"84820004",
		16#2045# => X"03ffff9f",
		16#2046# => X"e0845803",
		16#2047# => X"1000000c",
		16#2048# => X"bc470554",
		16#2049# => X"b8ee004f",
		16#204a# => X"9ce70077",
		16#204b# => X"03fffe5d",
		16#204c# => X"b8670003",
		16#204d# => X"85720004",
		16#204e# => X"e0a44008",
		16#204f# => X"a8830000",
		16#2050# => X"e0ab2804",
		16#2051# => X"03fffef5",
		16#2052# => X"d4122804",
		16#2053# => X"1000002a",
		16#2054# => X"15000000",
		16#2055# => X"b8ee0052",
		16#2056# => X"9ce7007c",
		16#2057# => X"03fffe51",
		16#2058# => X"b8670003",
		16#2059# => X"1000002c",
		16#205a# => X"bc430154",
		16#205b# => X"b904004c",
		16#205c# => X"03fffed5",
		16#205d# => X"9d08006e",
		16#205e# => X"9c600001",
		16#205f# => X"a8580000",
		16#2060# => X"d4181804",
		16#2061# => X"03ffff83",
		16#2062# => X"9c800000",
		16#2063# => X"a84c0000",
		16#2064# => X"a4a70003",
		16#2065# => X"bc250000",
		16#2066# => X"0c00003f",
		16#2067# => X"9c82fff8",
		16#2068# => X"84420000",
		16#2069# => X"e4222000",
		16#206a# => X"0ffffffa",
		16#206b# => X"9ce7ffff",
		16#206c# => X"e0631800",
		16#206d# => X"84520004",
		16#206e# => X"e4431000",
		16#206f# => X"13fffee2",
		16#2070# => X"bc030000",
		16#2071# => X"13fffee0",
		16#2072# => X"e0831003",
		16#2073# => X"bc240000",
		16#2074# => X"13fffe89",
		16#2075# => X"a8eb0000",
		16#2076# => X"e0631800",
		16#2077# => X"e0831003",
		16#2078# => X"bc040000",
		16#2079# => X"13fffffd",
		16#207a# => X"9d6b0004",
		16#207b# => X"03fffe82",
		16#207c# => X"a8eb0000",
		16#207d# => X"9c6003f0",
		16#207e# => X"03fffe2a",
		16#207f# => X"9ce0007e",
		16#2080# => X"84520008",
		16#2081# => X"9c60fffc",
		16#2082# => X"84820004",
		16#2083# => X"03ffff61",
		16#2084# => X"e0841803",
		16#2085# => X"1000001b",
		16#2086# => X"bc430554",
		16#2087# => X"b904004f",
		16#2088# => X"03fffea9",
		16#2089# => X"9d080077",
		16#208a# => X"a4a40fff",
		16#208b# => X"bc250000",
		16#208c# => X"13ffff15",
		16#208d# => X"15000000",
		16#208e# => X"e056a000",
		16#208f# => X"84920008",
		16#2090# => X"a8420001",
		16#2091# => X"03ffff42",
		16#2092# => X"d4041004",
		16#2093# => X"9c820008",
		16#2094# => X"18400001",
		16#2095# => X"a8700000",
		16#2096# => X"04001879",
		16#2097# => X"a8427a84",
		16#2098# => X"03ffff3b",
		16#2099# => X"84620000",
		16#209a# => X"03ffff21",
		16#209b# => X"9ec00000",
		16#209c# => X"18600001",
		16#209d# => X"a8636c14",
		16#209e# => X"03ffff09",
		16#209f# => X"d4035800",
		16#20a0# => X"13fffe91",
		16#20a1# => X"9d00007e",
		16#20a2# => X"b9040052",
		16#20a3# => X"03fffe8e",
		16#20a4# => X"9d08007c",
		16#20a5# => X"84920004",
		16#20a6# => X"ac43ffff",
		16#20a7# => X"e0441003",
		16#20a8# => X"03ffffc4",
		16#20a9# => X"d4121004",
		16#20aa# => X"44004800",
		16#20ab# => X"15000000",
		16#20ac# => X"44004800",
		16#20ad# => X"15000000",
		16#20ae# => X"b4600011",
		16#20af# => X"a8630020",
		16#20b0# => X"c0001840",
		16#20b1# => X"c0004820",
		16#20b2# => X"24000000",
		16#20b3# => X"15000000",
		16#20b4# => X"a8600020",
		16#20b5# => X"ac83ffff",
		16#20b6# => X"b4600011",
		16#20b7# => X"e0641803",
		16#20b8# => X"c0001840",
		16#20b9# => X"c0004820",
		16#20ba# => X"24000000",
		16#20bb# => X"15000000",
		16#20bc# => X"b4600011",
		16#20bd# => X"a8630040",
		16#20be# => X"c0001840",
		16#20bf# => X"c0004820",
		16#20c0# => X"24000000",
		16#20c1# => X"15000000",
		16#20c2# => X"a8600040",
		16#20c3# => X"ac83ffff",
		16#20c4# => X"b4600011",
		16#20c5# => X"e0641803",
		16#20c6# => X"c0001840",
		16#20c7# => X"c0004820",
		16#20c8# => X"24000000",
		16#20c9# => X"15000000",
		16#20ca# => X"b4600001",
		16#20cb# => X"a4830004",
		16#20cc# => X"e4040000",
		16#20cd# => X"10000021",
		16#20ce# => X"15000000",
		16#20cf# => X"b4c00011",
		16#20d0# => X"9ca0ffff",
		16#20d1# => X"aca50010",
		16#20d2# => X"e0a62803",
		16#20d3# => X"c0002811",
		16#20d4# => X"b4600006",
		16#20d5# => X"a4830080",
		16#20d6# => X"b8e40047",
		16#20d7# => X"a9000010",
		16#20d8# => X"e1c83808",
		16#20d9# => X"a4830078",
		16#20da# => X"b8e40043",
		16#20db# => X"a9000001",
		16#20dc# => X"e1a83808",
		16#20dd# => X"9cc00000",
		16#20de# => X"e0ae3808",
		16#20df# => X"c0803002",
		16#20e0# => X"e4262800",
		16#20e1# => X"13fffffe",
		16#20e2# => X"e0c67000",
		16#20e3# => X"b4c00011",
		16#20e4# => X"a8c60010",
		16#20e5# => X"c0003011",
		16#20e6# => X"15000000",
		16#20e7# => X"15000000",
		16#20e8# => X"15000000",
		16#20e9# => X"15000000",
		16#20ea# => X"15000000",
		16#20eb# => X"15000000",
		16#20ec# => X"15000000",
		16#20ed# => X"15000000",
		16#20ee# => X"b4600001",
		16#20ef# => X"a4830002",
		16#20f0# => X"e4040000",
		16#20f1# => X"10000019",
		16#20f2# => X"15000000",
		16#20f3# => X"b4c00011",
		16#20f4# => X"9ca0ffff",
		16#20f5# => X"aca50008",
		16#20f6# => X"e0a62803",
		16#20f7# => X"c0002811",
		16#20f8# => X"b4600005",
		16#20f9# => X"a4830080",
		16#20fa# => X"b8e40047",
		16#20fb# => X"a9000010",
		16#20fc# => X"e1c83808",
		16#20fd# => X"a4830078",
		16#20fe# => X"b8e40043",
		16#20ff# => X"a9000001",
		16#2100# => X"e1a83808",
		16#2101# => X"9cc00000",
		16#2102# => X"e0ae3808",
		16#2103# => X"c0603003",
		16#2104# => X"e4262800",
		16#2105# => X"13fffffe",
		16#2106# => X"e0c67000",
		16#2107# => X"b4c00011",
		16#2108# => X"a8c60008",
		16#2109# => X"c0003011",
		16#210a# => X"44004800",
		16#210b# => X"15000000",
		16#210c# => X"b5a00011",
		16#210d# => X"a9ad0010",
		16#210e# => X"c0006811",
		16#210f# => X"15000000",
		16#2110# => X"15000000",
		16#2111# => X"15000000",
		16#2112# => X"15000000",
		16#2113# => X"15000000",
		16#2114# => X"44004800",
		16#2115# => X"15000000",
		16#2116# => X"b5a00011",
		16#2117# => X"9d80ffff",
		16#2118# => X"ad8c0010",
		16#2119# => X"e18d6003",
		16#211a# => X"c0006011",
		16#211b# => X"44004800",
		16#211c# => X"15000000",
		16#211d# => X"44004800",
		16#211e# => X"c0801802",
		16#211f# => X"b5a00011",
		16#2120# => X"a9ad0008",
		16#2121# => X"c0006811",
		16#2122# => X"15000000",
		16#2123# => X"15000000",
		16#2124# => X"15000000",
		16#2125# => X"15000000",
		16#2126# => X"15000000",
		16#2127# => X"44004800",
		16#2128# => X"15000000",
		16#2129# => X"b5a00011",
		16#212a# => X"9d80ffff",
		16#212b# => X"ad8c0008",
		16#212c# => X"e18d6003",
		16#212d# => X"c0006011",
		16#212e# => X"44004800",
		16#212f# => X"15000000",
		16#2130# => X"44004800",
		16#2131# => X"c0601803",
		16#2132# => X"9c21fff4",
		16#2133# => X"d4014800",
		16#2134# => X"b4604802",
		16#2135# => X"18e00001",
		16#2136# => X"a8e76c18",
		16#2137# => X"1900ffff",
		16#2138# => X"a908ffff",
		16#2139# => X"19800001",
		16#213a# => X"a98c6c98",
		16#213b# => X"e083000f",
		16#213c# => X"e4240000",
		16#213d# => X"0c000014",
		16#213e# => X"15000000",
		16#213f# => X"9ca4ffff",
		16#2140# => X"b8c50002",
		16#2141# => X"e1c63800",
		16#2142# => X"e1a66000",
		16#2143# => X"85ce0000",
		16#2144# => X"e42e4000",
		16#2145# => X"0c000008",
		16#2146# => X"15000000",
		16#2147# => X"d4011804",
		16#2148# => X"846d0000",
		16#2149# => X"48007000",
		16#214a# => X"d4012808",
		16#214b# => X"84610004",
		16#214c# => X"84a10008",
		16#214d# => X"a8c00001",
		16#214e# => X"e0c62808",
		16#214f# => X"03ffffec",
		16#2150# => X"e0633005",
		16#2151# => X"85210000",
		16#2152# => X"c1201802",
		16#2153# => X"44004800",
		16#2154# => X"9c21000c",
		16#2155# => X"9c21fffc",
		16#2156# => X"d4013000",
		16#2157# => X"b8630002",
		16#2158# => X"18c00001",
		16#2159# => X"a8c66c18",
		16#215a# => X"e0c61800",
		16#215b# => X"d4062000",
		16#215c# => X"18c00001",
		16#215d# => X"a8c66c98",
		16#215e# => X"e0c61800",
		16#215f# => X"d4062800",
		16#2160# => X"84c10000",
		16#2161# => X"44004800",
		16#2162# => X"9c210004",
		16#2163# => X"9c21fffc",
		16#2164# => X"d4012000",
		16#2165# => X"a8800001",
		16#2166# => X"e0841808",
		16#2167# => X"b4604800",
		16#2168# => X"e0632004",
		16#2169# => X"c1201800",
		16#216a# => X"84810000",
		16#216b# => X"44004800",
		16#216c# => X"9c210004",
		16#216d# => X"9c21fffc",
		16#216e# => X"d4012000",
		16#216f# => X"a8800001",
		16#2170# => X"e0841808",
		16#2171# => X"ac84ffff",
		16#2172# => X"b4604800",
		16#2173# => X"e0632003",
		16#2174# => X"c1201800",
		16#2175# => X"84810000",
		16#2176# => X"44004800",
		16#2177# => X"9c210004",
		16#2178# => X"d4011000",
		16#2179# => X"d401280c",
		16#217a# => X"d4013010",
		16#217b# => X"d4013814",
		16#217c# => X"d4014018",
		16#217d# => X"d401481c",
		16#217e# => X"d4015020",
		16#217f# => X"d4015824",
		16#2180# => X"d4016028",
		16#2181# => X"d401682c",
		16#2182# => X"d4017030",
		16#2183# => X"d4017834",
		16#2184# => X"d4018038",
		16#2185# => X"d401883c",
		16#2186# => X"d4019040",
		16#2187# => X"d4019844",
		16#2188# => X"d401a048",
		16#2189# => X"d401a84c",
		16#218a# => X"d401b050",
		16#218b# => X"d401b854",
		16#218c# => X"d401c058",
		16#218d# => X"d401c85c",
		16#218e# => X"d401d060",
		16#218f# => X"d401d864",
		16#2190# => X"d401e068",
		16#2191# => X"d401e86c",
		16#2192# => X"d401f070",
		16#2193# => X"d401f874",
		16#2194# => X"a5a3ffff",
		16#2195# => X"b9ad0046",
		16#2196# => X"9dadfff8",
		16#2197# => X"19c00001",
		16#2198# => X"a9ce6d18",
		16#2199# => X"e1ce6800",
		16#219a# => X"85ae0000",
		16#219b# => X"19e0ffff",
		16#219c# => X"a9efffff",
		16#219d# => X"e42d7800",
		16#219e# => X"0c000025",
		16#219f# => X"15000000",
		16#21a0# => X"48006800",
		16#21a1# => X"e0642004",
		16#21a2# => X"84410000",
		16#21a3# => X"84610004",
		16#21a4# => X"84810008",
		16#21a5# => X"84a1000c",
		16#21a6# => X"84c10010",
		16#21a7# => X"84e10014",
		16#21a8# => X"85010018",
		16#21a9# => X"8521001c",
		16#21aa# => X"85410020",
		16#21ab# => X"85610024",
		16#21ac# => X"85810028",
		16#21ad# => X"85a1002c",
		16#21ae# => X"85c10030",
		16#21af# => X"85e10034",
		16#21b0# => X"86010038",
		16#21b1# => X"8621003c",
		16#21b2# => X"86410040",
		16#21b3# => X"86610044",
		16#21b4# => X"86810048",
		16#21b5# => X"86a1004c",
		16#21b6# => X"86c10050",
		16#21b7# => X"86e10054",
		16#21b8# => X"87010058",
		16#21b9# => X"8721005c",
		16#21ba# => X"87410060",
		16#21bb# => X"87610064",
		16#21bc# => X"87810068",
		16#21bd# => X"87a1006c",
		16#21be# => X"87c10070",
		16#21bf# => X"87e10074",
		16#21c0# => X"9c210100",
		16#21c1# => X"24000000",
		16#21c2# => X"15000000",
		16#21c3# => X"07fffc72",
		16#21c4# => X"e0642004",
		16#21c5# => X"9c21fffc",
		16#21c6# => X"d4012800",
		16#21c7# => X"b8630002",
		16#21c8# => X"9c63fff8",
		16#21c9# => X"18a00001",
		16#21ca# => X"a8a56d18",
		16#21cb# => X"e0a51800",
		16#21cc# => X"d4052000",
		16#21cd# => X"84a10000",
		16#21ce# => X"44004800",
		16#21cf# => X"9c210004",
		16#21d0# => X"18600001",
		16#21d1# => X"18800001",
		16#21d2# => X"a8639ac8",
		16#21d3# => X"d7e117fc",
		16#21d4# => X"a8849acc",
		16#21d5# => X"18400fff",
		16#21d6# => X"84a30000",
		16#21d7# => X"84840000",
		16#21d8# => X"a842ffff",
		16#21d9# => X"9ca50001",
		16#21da# => X"e0841003",
		16#21db# => X"18406000",
		16#21dc# => X"d4032800",
		16#21dd# => X"9c21fffc",
		16#21de# => X"e0841004",
		16#21df# => X"9c605000",
		16#21e0# => X"c0032000",
		16#21e1# => X"9c210004",
		16#21e2# => X"44004800",
		16#21e3# => X"8441fffc",
		16#21e4# => X"9c630000",
		16#21e5# => X"15000002",
		16#21e6# => X"44004800",
		16#21e7# => X"15000000",
		16#21e8# => X"c0032000",
		16#21e9# => X"44004800",
		16#21ea# => X"15000000",
		16#21eb# => X"b5630000",
		16#21ec# => X"44004800",
		16#21ed# => X"15000000",
		16#21ee# => X"18600001",
		16#21ef# => X"d7e117fc",
		16#21f0# => X"a8636d8c",
		16#21f1# => X"18800001",
		16#21f2# => X"84a30000",
		16#21f3# => X"1840d000",
		16#21f4# => X"a5650001",
		16#21f5# => X"a8847aac",
		16#21f6# => X"a8420001",
		16#21f7# => X"e1605802",
		16#21f8# => X"b8a50041",
		16#21f9# => X"84c40000",
		16#21fa# => X"e16b1003",
		16#21fb# => X"9cc60001",
		16#21fc# => X"e16b2805",
		16#21fd# => X"9c21fffc",
		16#21fe# => X"d4043000",
		16#21ff# => X"d4035800",
		16#2200# => X"9c210004",
		16#2201# => X"44004800",
		16#2202# => X"8441fffc",
		16#2203# => X"a8830000",
		16#2204# => X"18600001",
		16#2205# => X"d7e14ffc",
		16#2206# => X"a86338f8",
		16#2207# => X"d7e117f8",
		16#2208# => X"84630000",
		16#2209# => X"9c21fff8",
		16#220a# => X"07fff0b7",
		16#220b# => X"9c400000",
		16#220c# => X"18a00001",
		16#220d# => X"18800000",
		16#220e# => X"a8a59acc",
		16#220f# => X"9c600005",
		16#2210# => X"d4055800",
		16#2211# => X"18a00001",
		16#2212# => X"a8848740",
		16#2213# => X"a8a59ac8",
		16#2214# => X"d4051000",
		16#2215# => X"9c210008",
		16#2216# => X"8521fffc",
		16#2217# => X"03ffffae",
		16#2218# => X"8441fff8",
		16#2219# => X"18600001",
		16#221a# => X"d7e117fc",
		16#221b# => X"a8639acc",
		16#221c# => X"18400fff",
		16#221d# => X"84830000",
		16#221e# => X"a842ffff",
		16#221f# => X"9c21fffc",
		16#2220# => X"e0841003",
		16#2221# => X"18406000",
		16#2222# => X"9c605000",
		16#2223# => X"e0841004",
		16#2224# => X"c0032000",
		16#2225# => X"9c600011",
		16#2226# => X"b4830000",
		16#2227# => X"a8840002",
		16#2228# => X"c0032000",
		16#2229# => X"9c210004",
		16#222a# => X"44004800",
		16#222b# => X"8441fffc",
		16#222c# => X"d7e117fc",
		16#222d# => X"9c600011",
		16#222e# => X"9c21fffc",
		16#222f# => X"b4830000",
		16#2230# => X"9c40fffd",
		16#2231# => X"e0841003",
		16#2232# => X"c0032000",
		16#2233# => X"9c210004",
		16#2234# => X"44004800",
		16#2235# => X"8441fffc",
		16#2236# => X"18600001",
		16#2237# => X"a8639ac8",
		16#2238# => X"85630000",
		16#2239# => X"44004800",
		16#223a# => X"15000000",
		16#223b# => X"18600001",
		16#223c# => X"d7e117fc",
		16#223d# => X"a8639ac8",
		16#223e# => X"9c400000",
		16#223f# => X"9c21fffc",
		16#2240# => X"d4031000",
		16#2241# => X"9c210004",
		16#2242# => X"44004800",
		16#2243# => X"8441fffc",
		16#2244# => X"d7e14ffc",
		16#2245# => X"9c21fffc",
		16#2246# => X"a8a40000",
		16#2247# => X"9cc10004",
		16#2248# => X"04000353",
		16#2249# => X"84830008",
		16#224a# => X"9c210004",
		16#224b# => X"8521fffc",
		16#224c# => X"44004800",
		16#224d# => X"15000000",
		16#224e# => X"a8a30000",
		16#224f# => X"18600001",
		16#2250# => X"d7e14ffc",
		16#2251# => X"a86363e0",
		16#2252# => X"9c21fffc",
		16#2253# => X"84630000",
		16#2254# => X"9cc10004",
		16#2255# => X"04000346",
		16#2256# => X"84830008",
		16#2257# => X"9c210004",
		16#2258# => X"8521fffc",
		16#2259# => X"44004800",
		16#225a# => X"15000000",
		16#225b# => X"d7e117f4",
		16#225c# => X"d7e177f8",
		16#225d# => X"d7e14ffc",
		16#225e# => X"a8430000",
		16#225f# => X"9c21ffd8",
		16#2260# => X"a8640000",
		16#2261# => X"040002fc",
		16#2262# => X"a9c40000",
		16#2263# => X"18600001",
		16#2264# => X"18e00001",
		16#2265# => X"a86363e0",
		16#2266# => X"9ccb0001",
		16#2267# => X"84630000",
		16#2268# => X"a8e73b53",
		16#2269# => X"84a30008",
		16#226a# => X"d4013808",
		16#226b# => X"9865000c",
		16#226c# => X"9ce00001",
		16#226d# => X"d4013018",
		16#226e# => X"9cc00002",
		16#226f# => X"a4832000",
		16#2270# => X"d4017000",
		16#2271# => X"d4015804",
		16#2272# => X"d401380c",
		16#2273# => X"d4010810",
		16#2274# => X"bc240000",
		16#2275# => X"10000008",
		16#2276# => X"d4013014",
		16#2277# => X"84850064",
		16#2278# => X"9cc0dfff",
		16#2279# => X"a8632000",
		16#227a# => X"e0843003",
		16#227b# => X"dc05180c",
		16#227c# => X"d4052064",
		16#227d# => X"a8620000",
		16#227e# => X"9ca10010",
		16#227f# => X"0400175c",
		16#2280# => X"84820008",
		16#2281# => X"bc0b0000",
		16#2282# => X"0c000008",
		16#2283# => X"9c60000a",
		16#2284# => X"9c210028",
		16#2285# => X"a9630000",
		16#2286# => X"8521fffc",
		16#2287# => X"8441fff4",
		16#2288# => X"44004800",
		16#2289# => X"85c1fff8",
		16#228a# => X"9c210028",
		16#228b# => X"9c60ffff",
		16#228c# => X"8521fffc",
		16#228d# => X"a9630000",
		16#228e# => X"8441fff4",
		16#228f# => X"44004800",
		16#2290# => X"85c1fff8",
		16#2291# => X"a8830000",
		16#2292# => X"18600001",
		16#2293# => X"d7e14ffc",
		16#2294# => X"a86363e0",
		16#2295# => X"9c21fffc",
		16#2296# => X"84630000",
		16#2297# => X"9c210004",
		16#2298# => X"8521fffc",
		16#2299# => X"03ffffc2",
		16#229a# => X"15000000",
		16#229b# => X"d7e197e0",
		16#229c# => X"aa430000",
		16#229d# => X"ac650004",
		16#229e# => X"d7e117d4",
		16#229f# => X"d7e1d7f0",
		16#22a0# => X"e0452800",
		16#22a1# => X"ab450000",
		16#22a2# => X"e0a01802",
		16#22a3# => X"e042d000",
		16#22a4# => X"e0651804",
		16#22a5# => X"b8ba0042",
		16#22a6# => X"b863005f",
		16#22a7# => X"d7e1a7e4",
		16#22a8# => X"d7e1b7e8",
		16#22a9# => X"d7e14ffc",
		16#22aa# => X"d7e177d8",
		16#22ab# => X"d7e187dc",
		16#22ac# => X"d7e1c7ec",
		16#22ad# => X"d7e1e7f4",
		16#22ae# => X"d7e1f7f8",
		16#22af# => X"aa860000",
		16#22b0# => X"9c21ffb0",
		16#22b1# => X"a4da0003",
		16#22b2# => X"e0421000",
		16#22b3# => X"d4012804",
		16#22b4# => X"d4011820",
		16#22b5# => X"d4012000",
		16#22b6# => X"d4013010",
		16#22b7# => X"d4011014",
		16#22b8# => X"e2c0d002",
		16#22b9# => X"a4520003",
		16#22ba# => X"bc220000",
		16#22bb# => X"10000007",
		16#22bc# => X"9f000002",
		16#22bd# => X"84e10010",
		16#22be# => X"bc270000",
		16#22bf# => X"10000004",
		16#22c0# => X"84410000",
		16#22c1# => X"87010020",
		16#22c2# => X"84410000",
		16#22c3# => X"bc420006",
		16#22c4# => X"0c0001fe",
		16#22c5# => X"84610000",
		16#22c6# => X"abd20000",
		16#22c7# => X"b8430041",
		16#22c8# => X"bc230007",
		16#22c9# => X"e042d306",
		16#22ca# => X"100000ba",
		16#22cb# => X"e0521000",
		16#22cc# => X"84810014",
		16#22cd# => X"e1d22000",
		16#22ce# => X"bc380000",
		16#22cf# => X"100000d1",
		16#22d0# => X"e0f2d000",
		16#22d1# => X"84820000",
		16#22d2# => X"84720000",
		16#22d3# => X"d4122000",
		16#22d4# => X"d4021800",
		16#22d5# => X"a84e0000",
		16#22d6# => X"d401380c",
		16#22d7# => X"aa070000",
		16#22d8# => X"d4013808",
		16#22d9# => X"9f800000",
		16#22da# => X"e4501000",
		16#22db# => X"0c00003b",
		16#22dc# => X"a8700000",
		16#22dd# => X"bc3c0000",
		16#22de# => X"0c00019c",
		16#22df# => X"84610000",
		16#22e0# => X"84810008",
		16#22e1# => X"e383d306",
		16#22e2# => X"e0a49002",
		16#22e3# => X"e0702002",
		16#22e4# => X"e5a51800",
		16#22e5# => X"10000003",
		16#22e6# => X"e392e000",
		16#22e7# => X"a8a30000",
		16#22e8# => X"bda50000",
		16#22e9# => X"1000000d",
		16#22ea# => X"bc180002",
		16#22eb# => X"e0902802",
		16#22ec# => X"0c000103",
		16#22ed# => X"e0d22800",
		16#22ee# => X"8ce40000",
		16#22ef# => X"90be0000",
		16#22f0# => X"d81e3800",
		16#22f1# => X"d8042800",
		16#22f2# => X"9fde0001",
		16#22f3# => X"e43e3000",
		16#22f4# => X"13fffffa",
		16#22f5# => X"9c840001",
		16#22f6# => X"e0dc7002",
		16#22f7# => X"e04e1002",
		16#22f8# => X"e0c6d002",
		16#22f9# => X"e4a61000",
		16#22fa# => X"10000004",
		16#22fb# => X"bda60000",
		16#22fc# => X"a8c20000",
		16#22fd# => X"bda60000",
		16#22fe# => X"1000000e",
		16#22ff# => X"a8a60000",
		16#2300# => X"bc180002",
		16#2301# => X"0c0000e2",
		16#2302# => X"e09c3002",
		16#2303# => X"8ce40000",
		16#2304# => X"90d00000",
		16#2305# => X"d8103800",
		16#2306# => X"d8043000",
		16#2307# => X"9ca5ffff",
		16#2308# => X"9e100001",
		16#2309# => X"bc250000",
		16#230a# => X"13fffff9",
		16#230b# => X"9c840001",
		16#230c# => X"e47a1800",
		16#230d# => X"0c0000a2",
		16#230e# => X"e47a1000",
		16#230f# => X"100000aa",
		16#2310# => X"a8620000",
		16#2311# => X"a89a0000",
		16#2312# => X"07ffefaf",
		16#2313# => X"e25c1002",
		16#2314# => X"03ffffa5",
		16#2315# => X"d4015800",
		16#2316# => X"4800a000",
		16#2317# => X"a8920000",
		16#2318# => X"bdab0000",
		16#2319# => X"0c00000e",
		16#231a# => X"a8620000",
		16#231b# => X"0000004e",
		16#231c# => X"bc2b0000",
		16#231d# => X"84ae0000",
		16#231e# => X"84620000",
		16#231f# => X"d4022800",
		16#2320# => X"d40e1800",
		16#2321# => X"e1ceb000",
		16#2322# => X"9f800001",
		16#2323# => X"e042b000",
		16#2324# => X"e4b01000",
		16#2325# => X"0fffffb8",
		16#2326# => X"a8620000",
		16#2327# => X"4800a000",
		16#2328# => X"a8920000",
		16#2329# => X"bd6b0000",
		16#232a# => X"0c000015",
		16#232b# => X"bc0b0000",
		16#232c# => X"0ffffff7",
		16#232d# => X"bc380000",
		16#232e# => X"0fffffef",
		16#232f# => X"bc380001",
		16#2330# => X"0c00001d",
		16#2331# => X"a90e0000",
		16#2332# => X"a87a0000",
		16#2333# => X"a8e20000",
		16#2334# => X"8c880000",
		16#2335# => X"90c70000",
		16#2336# => X"d8072000",
		16#2337# => X"d8083000",
		16#2338# => X"9c63ffff",
		16#2339# => X"9ce70001",
		16#233a# => X"bd430000",
		16#233b# => X"13fffff9",
		16#233c# => X"9d080001",
		16#233d# => X"03ffffe5",
		16#233e# => X"e1ceb000",
		16#233f# => X"e4501000",
		16#2340# => X"13ffff9d",
		16#2341# => X"a8c20000",
		16#2342# => X"bc380000",
		16#2343# => X"10000018",
		16#2344# => X"bc380001",
		16#2345# => X"84620000",
		16#2346# => X"84500000",
		16#2347# => X"d4101800",
		16#2348# => X"d4061000",
		16#2349# => X"e210d000",
		16#234a# => X"e046b000",
		16#234b# => X"03ffff8f",
		16#234c# => X"9f800001",
		16#234d# => X"a8c20000",
		16#234e# => X"a86e0000",
		16#234f# => X"84e10004",
		16#2350# => X"85030000",
		16#2351# => X"84a60000",
		16#2352# => X"d4064000",
		16#2353# => X"d4032800",
		16#2354# => X"9ce7ffff",
		16#2355# => X"9cc60004",
		16#2356# => X"bd470000",
		16#2357# => X"13fffff9",
		16#2358# => X"9c630004",
		16#2359# => X"03ffffc9",
		16#235a# => X"e1ceb000",
		16#235b# => X"0c00001c",
		16#235c# => X"a8ba0000",
		16#235d# => X"a8700000",
		16#235e# => X"8c820000",
		16#235f# => X"90e30000",
		16#2360# => X"d8032000",
		16#2361# => X"d8023800",
		16#2362# => X"9ca5ffff",
		16#2363# => X"9c630001",
		16#2364# => X"bd450000",
		16#2365# => X"13fffff9",
		16#2366# => X"9c420001",
		16#2367# => X"03ffffe3",
		16#2368# => X"e210d000",
		16#2369# => X"1000000c",
		16#236a# => X"bc380000",
		16#236b# => X"1000005b",
		16#236c# => X"84a10008",
		16#236d# => X"84900000",
		16#236e# => X"84650000",
		16#236f# => X"d4052000",
		16#2370# => X"d4101800",
		16#2371# => X"84610008",
		16#2372# => X"9f800001",
		16#2373# => X"e063d000",
		16#2374# => X"d4011808",
		16#2375# => X"03ffff65",
		16#2376# => X"e210d000",
		16#2377# => X"a8700000",
		16#2378# => X"84a10004",
		16#2379# => X"84e20000",
		16#237a# => X"84830000",
		16#237b# => X"d4033800",
		16#237c# => X"d4022000",
		16#237d# => X"9ca5ffff",
		16#237e# => X"9c630004",
		16#237f# => X"bd450000",
		16#2380# => X"13fffff9",
		16#2381# => X"9c420004",
		16#2382# => X"03ffffc8",
		16#2383# => X"e210d000",
		16#2384# => X"84a10000",
		16#2385# => X"9dc5ffff",
		16#2386# => X"bca50028",
		16#2387# => X"e1ced306",
		16#2388# => X"0c000074",
		16#2389# => X"e1d27000",
		16#238a# => X"ab8e0000",
		16#238b# => X"aa120000",
		16#238c# => X"a8700000",
		16#238d# => X"4800a000",
		16#238e# => X"a8820000",
		16#238f# => X"bd6b0000",
		16#2390# => X"0c000046",
		16#2391# => X"a8620000",
		16#2392# => X"4800a000",
		16#2393# => X"a89c0000",
		16#2394# => X"bd4b0000",
		16#2395# => X"13ffff3a",
		16#2396# => X"bc380000",
		16#2397# => X"a8700000",
		16#2398# => X"a89c0000",
		16#2399# => X"4800a000",
		16#239a# => X"a85c0000",
		16#239b# => X"bd6b0000",
		16#239c# => X"13ffff33",
		16#239d# => X"bc380000",
		16#239e# => X"03ffff31",
		16#239f# => X"a8500000",
		16#23a0# => X"bc380001",
		16#23a1# => X"0c000097",
		16#23a2# => X"a8ba0000",
		16#23a3# => X"a8720000",
		16#23a4# => X"8cc20000",
		16#23a5# => X"90830000",
		16#23a6# => X"d8033000",
		16#23a7# => X"d8022000",
		16#23a8# => X"9ca5ffff",
		16#23a9# => X"9c630001",
		16#23aa# => X"bd450000",
		16#23ab# => X"13fffff9",
		16#23ac# => X"9c420001",
		16#23ad# => X"03ffff28",
		16#23ae# => X"e0f2d000",
		16#23af# => X"07ffef12",
		16#23b0# => X"a89a0000",
		16#23b1# => X"a8720000",
		16#23b2# => X"a88b0000",
		16#23b3# => X"a8ba0000",
		16#23b4# => X"07fffee7",
		16#23b5# => X"a8d40000",
		16#23b6# => X"e47a1000",
		16#23b7# => X"0fffff5a",
		16#23b8# => X"a8620000",
		16#23b9# => X"9c210050",
		16#23ba# => X"8521fffc",
		16#23bb# => X"8441ffd4",
		16#23bc# => X"85c1ffd8",
		16#23bd# => X"8601ffdc",
		16#23be# => X"8641ffe0",
		16#23bf# => X"8681ffe4",
		16#23c0# => X"86c1ffe8",
		16#23c1# => X"8701ffec",
		16#23c2# => X"8741fff0",
		16#23c3# => X"8781fff4",
		16#23c4# => X"44004800",
		16#23c5# => X"87c1fff8",
		16#23c6# => X"bc380001",
		16#23c7# => X"0c00007e",
		16#23c8# => X"a8ba0000",
		16#23c9# => X"a8900000",
		16#23ca# => X"84610008",
		16#23cb# => X"8ce40000",
		16#23cc# => X"90c30000",
		16#23cd# => X"d8033800",
		16#23ce# => X"d8043000",
		16#23cf# => X"9ca5ffff",
		16#23d0# => X"9c630001",
		16#23d1# => X"bd450000",
		16#23d2# => X"13fffff9",
		16#23d3# => X"9c840001",
		16#23d4# => X"03ffff9e",
		16#23d5# => X"84610008",
		16#23d6# => X"4800a000",
		16#23d7# => X"a89c0000",
		16#23d8# => X"bd8b0000",
		16#23d9# => X"13fffef5",
		16#23da# => X"a8700000",
		16#23db# => X"a89c0000",
		16#23dc# => X"4800a000",
		16#23dd# => X"a8500000",
		16#23de# => X"bd6b0000",
		16#23df# => X"13fffef0",
		16#23e0# => X"bc380000",
		16#23e1# => X"03fffeee",
		16#23e2# => X"a85c0000",
		16#23e3# => X"b8c60042",
		16#23e4# => X"84e40000",
		16#23e5# => X"84b00000",
		16#23e6# => X"d4103800",
		16#23e7# => X"d4042800",
		16#23e8# => X"9cc6ffff",
		16#23e9# => X"9e100004",
		16#23ea# => X"bd460000",
		16#23eb# => X"13fffff9",
		16#23ec# => X"9c840004",
		16#23ed# => X"03ffff20",
		16#23ee# => X"e47a1800",
		16#23ef# => X"b8a50042",
		16#23f0# => X"a8d20000",
		16#23f1# => X"85040000",
		16#23f2# => X"84e60000",
		16#23f3# => X"d4064000",
		16#23f4# => X"d4043800",
		16#23f5# => X"9ca5ffff",
		16#23f6# => X"9cc60004",
		16#23f7# => X"bd450000",
		16#23f8# => X"13fffff9",
		16#23f9# => X"9c840004",
		16#23fa# => X"03fffefd",
		16#23fb# => X"e0dc7002",
		16#23fc# => X"b8850043",
		16#23fd# => X"a8720000",
		16#23fe# => X"e084d306",
		16#23ff# => X"e0c42000",
		16#2400# => X"e2122000",
		16#2401# => X"d4012008",
		16#2402# => X"d401301c",
		16#2403# => X"a8900000",
		16#2404# => X"4800a000",
		16#2405# => X"e3923000",
		16#2406# => X"bd6b0000",
		16#2407# => X"0c000066",
		16#2408# => X"a8700000",
		16#2409# => X"4800a000",
		16#240a# => X"a89c0000",
		16#240b# => X"bd4b0000",
		16#240c# => X"0c000105",
		16#240d# => X"a8720000",
		16#240e# => X"84e10008",
		16#240f# => X"84a10008",
		16#2410# => X"e0e03802",
		16#2411# => X"a8820000",
		16#2412# => X"e0623800",
		16#2413# => X"d4013818",
		16#2414# => X"d401180c",
		16#2415# => X"4800a000",
		16#2416# => X"e3822800",
		16#2417# => X"bd6b0000",
		16#2418# => X"0c000048",
		16#2419# => X"a8620000",
		16#241a# => X"4800a000",
		16#241b# => X"a89c0000",
		16#241c# => X"bd4b0000",
		16#241d# => X"0c0000ec",
		16#241e# => X"8461000c",
		16#241f# => X"84c1001c",
		16#2420# => X"84e10018",
		16#2421# => X"e0ce3002",
		16#2422# => X"e38e3800",
		16#2423# => X"d4013008",
		16#2424# => X"a8660000",
		16#2425# => X"4800a000",
		16#2426# => X"a89c0000",
		16#2427# => X"bd6b0000",
		16#2428# => X"0c00002b",
		16#2429# => X"a87c0000",
		16#242a# => X"4800a000",
		16#242b# => X"a88e0000",
		16#242c# => X"bd4b0000",
		16#242d# => X"13ffff60",
		16#242e# => X"a8700000",
		16#242f# => X"84610008",
		16#2430# => X"a88e0000",
		16#2431# => X"4800a000",
		16#2432# => X"ab8e0000",
		16#2433# => X"bd6b0000",
		16#2434# => X"13ffff59",
		16#2435# => X"a8700000",
		16#2436# => X"03ffff57",
		16#2437# => X"87810008",
		16#2438# => X"a8720000",
		16#2439# => X"84810004",
		16#243a# => X"84c20000",
		16#243b# => X"84a30000",
		16#243c# => X"d4033000",
		16#243d# => X"d4022800",
		16#243e# => X"9c84ffff",
		16#243f# => X"9c630004",
		16#2440# => X"bd440000",
		16#2441# => X"13fffff9",
		16#2442# => X"9c420004",
		16#2443# => X"03fffe92",
		16#2444# => X"e0f2d000",
		16#2445# => X"84810008",
		16#2446# => X"a8700000",
		16#2447# => X"84a10004",
		16#2448# => X"84e30000",
		16#2449# => X"84c40000",
		16#244a# => X"d4043800",
		16#244b# => X"d4033000",
		16#244c# => X"9ca5ffff",
		16#244d# => X"9c840004",
		16#244e# => X"bd450000",
		16#244f# => X"13fffff9",
		16#2450# => X"9c630004",
		16#2451# => X"03ffff21",
		16#2452# => X"84610008",
		16#2453# => X"4800a000",
		16#2454# => X"a88e0000",
		16#2455# => X"bd8b0000",
		16#2456# => X"13ffff36",
		16#2457# => X"84610008",
		16#2458# => X"a88e0000",
		16#2459# => X"4800a000",
		16#245a# => X"ab830000",
		16#245b# => X"bd6b0000",
		16#245c# => X"13ffff31",
		16#245d# => X"a8700000",
		16#245e# => X"03ffff2f",
		16#245f# => X"ab8e0000",
		16#2460# => X"4800a000",
		16#2461# => X"a89c0000",
		16#2462# => X"bd8b0000",
		16#2463# => X"13ffffbc",
		16#2464# => X"8461000c",
		16#2465# => X"a89c0000",
		16#2466# => X"4800a000",
		16#2467# => X"a8430000",
		16#2468# => X"bd6b0000",
		16#2469# => X"13ffffb7",
		16#246a# => X"84c1001c",
		16#246b# => X"03ffffb5",
		16#246c# => X"a85c0000",
		16#246d# => X"4800a000",
		16#246e# => X"a89c0000",
		16#246f# => X"bd8b0000",
		16#2470# => X"13ffff9e",
		16#2471# => X"a8720000",
		16#2472# => X"a89c0000",
		16#2473# => X"4800a000",
		16#2474# => X"aa120000",
		16#2475# => X"bd6b0000",
		16#2476# => X"13ffff99",
		16#2477# => X"84e10008",
		16#2478# => X"03ffff97",
		16#2479# => X"aa1c0000",
		16#247a# => X"84a10000",
		16#247b# => X"84c1000c",
		16#247c# => X"e045d306",
		16#247d# => X"e0521000",
		16#247e# => X"e4a23000",
		16#247f# => X"13ffff3a",
		16#2480# => X"d4011000",
		16#2481# => X"e2c0d002",
		16#2482# => X"ab860000",
		16#2483# => X"e3c6b000",
		16#2484# => X"e472e000",
		16#2485# => X"10000028",
		16#2486# => X"a85c0000",
		16#2487# => X"0000000c",
		16#2488# => X"a9de0000",
		16#2489# => X"e050b002",
		16#248a# => X"848e0000",
		16#248b# => X"84620000",
		16#248c# => X"d4022000",
		16#248d# => X"d40e1800",
		16#248e# => X"e1ceb000",
		16#248f# => X"e04eb002",
		16#2490# => X"e4721000",
		16#2491# => X"1000001c",
		16#2492# => X"a8500000",
		16#2493# => X"e202b000",
		16#2494# => X"a8820000",
		16#2495# => X"4800a000",
		16#2496# => X"a8700000",
		16#2497# => X"bd4b0000",
		16#2498# => X"0c000015",
		16#2499# => X"bc380000",
		16#249a# => X"0fffffef",
		16#249b# => X"bc380001",
		16#249c# => X"0c000018",
		16#249d# => X"a8ba0000",
		16#249e# => X"a8900000",
		16#249f# => X"8ce40000",
		16#24a0# => X"90620000",
		16#24a1# => X"d8023800",
		16#24a2# => X"d8041800",
		16#24a3# => X"9ca5ffff",
		16#24a4# => X"9c420001",
		16#24a5# => X"bd450000",
		16#24a6# => X"13fffff9",
		16#24a7# => X"9c840001",
		16#24a8# => X"e1ceb000",
		16#24a9# => X"e04eb002",
		16#24aa# => X"e4721000",
		16#24ab# => X"0fffffe8",
		16#24ac# => X"a8500000",
		16#24ad# => X"e39cd000",
		16#24ae# => X"84410000",
		16#24af# => X"e4a2e000",
		16#24b0# => X"0fffffd4",
		16#24b1# => X"e3ded000",
		16#24b2# => X"03ffff08",
		16#24b3# => X"9c210050",
		16#24b4# => X"e070b002",
		16#24b5# => X"a84e0000",
		16#24b6# => X"84810004",
		16#24b7# => X"84c20000",
		16#24b8# => X"84a30000",
		16#24b9# => X"d4033000",
		16#24ba# => X"d4022800",
		16#24bb# => X"9c84ffff",
		16#24bc# => X"9c630004",
		16#24bd# => X"bd440000",
		16#24be# => X"13fffff9",
		16#24bf# => X"9c420004",
		16#24c0# => X"03ffffcf",
		16#24c1# => X"e1ceb000",
		16#24c2# => X"e042d306",
		16#24c3# => X"e0521000",
		16#24c4# => X"e3d2d000",
		16#24c5# => X"e47e1000",
		16#24c6# => X"13fffef3",
		16#24c7# => X"d4011000",
		16#24c8# => X"e2c0d002",
		16#24c9# => X"ab9e0000",
		16#24ca# => X"e3deb000",
		16#24cb# => X"e472e000",
		16#24cc# => X"10000028",
		16#24cd# => X"a85c0000",
		16#24ce# => X"0000000c",
		16#24cf# => X"a9de0000",
		16#24d0# => X"e050b002",
		16#24d1# => X"848e0000",
		16#24d2# => X"84620000",
		16#24d3# => X"d4022000",
		16#24d4# => X"d40e1800",
		16#24d5# => X"e1ceb000",
		16#24d6# => X"e04eb002",
		16#24d7# => X"e4721000",
		16#24d8# => X"1000001c",
		16#24d9# => X"a8500000",
		16#24da# => X"e202b000",
		16#24db# => X"a8820000",
		16#24dc# => X"4800a000",
		16#24dd# => X"a8700000",
		16#24de# => X"bd4b0000",
		16#24df# => X"0c000015",
		16#24e0# => X"bc380000",
		16#24e1# => X"0fffffef",
		16#24e2# => X"bc380001",
		16#24e3# => X"0c000018",
		16#24e4# => X"a8ba0000",
		16#24e5# => X"a8900000",
		16#24e6# => X"8cc40000",
		16#24e7# => X"90620000",
		16#24e8# => X"d8023000",
		16#24e9# => X"d8041800",
		16#24ea# => X"9ca5ffff",
		16#24eb# => X"9c420001",
		16#24ec# => X"bd450000",
		16#24ed# => X"13fffff9",
		16#24ee# => X"9c840001",
		16#24ef# => X"e1ceb000",
		16#24f0# => X"e04eb002",
		16#24f1# => X"e4721000",
		16#24f2# => X"0fffffe8",
		16#24f3# => X"a8500000",
		16#24f4# => X"e39cd000",
		16#24f5# => X"84e10000",
		16#24f6# => X"e47c3800",
		16#24f7# => X"0fffffd4",
		16#24f8# => X"e3ded000",
		16#24f9# => X"03fffec1",
		16#24fa# => X"9c210050",
		16#24fb# => X"e070b002",
		16#24fc# => X"a84e0000",
		16#24fd# => X"84810004",
		16#24fe# => X"84c20000",
		16#24ff# => X"84a30000",
		16#2500# => X"d4033000",
		16#2501# => X"d4022800",
		16#2502# => X"9c84ffff",
		16#2503# => X"9c630004",
		16#2504# => X"bd440000",
		16#2505# => X"13fffff9",
		16#2506# => X"9c420004",
		16#2507# => X"03ffffcf",
		16#2508# => X"e1ceb000",
		16#2509# => X"a89c0000",
		16#250a# => X"4800a000",
		16#250b# => X"a85c0000",
		16#250c# => X"bd6b0000",
		16#250d# => X"13ffff13",
		16#250e# => X"84c1001c",
		16#250f# => X"03ffff11",
		16#2510# => X"8441000c",
		16#2511# => X"a89c0000",
		16#2512# => X"4800a000",
		16#2513# => X"aa1c0000",
		16#2514# => X"bd6b0000",
		16#2515# => X"13fffefa",
		16#2516# => X"84e10008",
		16#2517# => X"03fffef8",
		16#2518# => X"aa120000",
		16#2519# => X"18800001",
		16#251a# => X"d7e117fc",
		16#251b# => X"a88463e0",
		16#251c# => X"9c400000",
		16#251d# => X"84840000",
		16#251e# => X"9c21fffc",
		16#251f# => X"d40418a8",
		16#2520# => X"d40410a4",
		16#2521# => X"9c210004",
		16#2522# => X"44004800",
		16#2523# => X"8441fffc",
		16#2524# => X"d7e117f8",
		16#2525# => X"18400001",
		16#2526# => X"18a05851",
		16#2527# => X"18c04c95",
		16#2528# => X"a84263e0",
		16#2529# => X"d7e14ffc",
		16#252a# => X"a8a5f42d",
		16#252b# => X"9c21fff8",
		16#252c# => X"84420000",
		16#252d# => X"846200a4",
		16#252e# => X"848200a8",
		16#252f# => X"07fff898",
		16#2530# => X"a8c67f2d",
		16#2531# => X"9c600001",
		16#2532# => X"bc6cffff",
		16#2533# => X"10000003",
		16#2534# => X"9c8c0001",
		16#2535# => X"9c600000",
		16#2536# => X"e1635800",
		16#2537# => X"d40220a8",
		16#2538# => X"d40258a4",
		16#2539# => X"9c210008",
		16#253a# => X"18407fff",
		16#253b# => X"8521fffc",
		16#253c# => X"a842ffff",
		16#253d# => X"e16b1003",
		16#253e# => X"44004800",
		16#253f# => X"8441fff8",
		16#2540# => X"d7e117f4",
		16#2541# => X"18400001",
		16#2542# => X"d7e177f8",
		16#2543# => X"a8429ad0",
		16#2544# => X"a9c30000",
		16#2545# => X"a8640000",
		16#2546# => X"9c800000",
		16#2547# => X"d7e14ffc",
		16#2548# => X"d4022000",
		16#2549# => X"04002853",
		16#254a# => X"9c21fff4",
		16#254b# => X"bc2bffff",
		16#254c# => X"0c000007",
		16#254d# => X"15000000",
		16#254e# => X"9c21000c",
		16#254f# => X"8521fffc",
		16#2550# => X"8441fff4",
		16#2551# => X"44004800",
		16#2552# => X"85c1fff8",
		16#2553# => X"84420000",
		16#2554# => X"bc020000",
		16#2555# => X"13fffff9",
		16#2556# => X"15000000",
		16#2557# => X"d40e1000",
		16#2558# => X"9c21000c",
		16#2559# => X"8521fffc",
		16#255a# => X"8441fff4",
		16#255b# => X"44004800",
		16#255c# => X"85c1fff8",
		16#255d# => X"d7e117fc",
		16#255e# => X"a4830003",
		16#255f# => X"bc040000",
		16#2560# => X"10000039",
		16#2561# => X"9c21fffc",
		16#2562# => X"91630000",
		16#2563# => X"bc0b0000",
		16#2564# => X"10000032",
		16#2565# => X"15000000",
		16#2566# => X"00000006",
		16#2567# => X"a9630000",
		16#2568# => X"908b0000",
		16#2569# => X"bc240000",
		16#256a# => X"0c00002b",
		16#256b# => X"15000000",
		16#256c# => X"9d6b0001",
		16#256d# => X"a48b0003",
		16#256e# => X"bc240000",
		16#256f# => X"13fffff9",
		16#2570# => X"15000000",
		16#2571# => X"1840fefe",
		16#2572# => X"848b0000",
		16#2573# => X"a842feff",
		16#2574# => X"e0a41000",
		16#2575# => X"ac84ffff",
		16#2576# => X"18408080",
		16#2577# => X"e0852003",
		16#2578# => X"a8428080",
		16#2579# => X"e0841003",
		16#257a# => X"bc240000",
		16#257b# => X"10000010",
		16#257c# => X"15000000",
		16#257d# => X"9d6b0004",
		16#257e# => X"1840fefe",
		16#257f# => X"848b0000",
		16#2580# => X"a842feff",
		16#2581# => X"e0a41000",
		16#2582# => X"ac84ffff",
		16#2583# => X"18408080",
		16#2584# => X"e0852003",
		16#2585# => X"a8428080",
		16#2586# => X"e0841003",
		16#2587# => X"bc040000",
		16#2588# => X"13fffff6",
		16#2589# => X"9d6b0004",
		16#258a# => X"9d6bfffc",
		16#258b# => X"908b0000",
		16#258c# => X"bc040000",
		16#258d# => X"10000008",
		16#258e# => X"15000000",
		16#258f# => X"9d6b0001",
		16#2590# => X"908b0000",
		16#2591# => X"bc240000",
		16#2592# => X"13fffffe",
		16#2593# => X"9d6b0001",
		16#2594# => X"9d6bffff",
		16#2595# => X"e16b1802",
		16#2596# => X"9c210004",
		16#2597# => X"44004800",
		16#2598# => X"8441fffc",
		16#2599# => X"03ffffd8",
		16#259a# => X"a9630000",
		16#259b# => X"d7e14ffc",
		16#259c# => X"d7e117d4",
		16#259d# => X"d7e177d8",
		16#259e# => X"d7e187dc",
		16#259f# => X"d7e197e0",
		16#25a0# => X"d7e1a7e4",
		16#25a1# => X"d7e1b7e8",
		16#25a2# => X"d7e1c7ec",
		16#25a3# => X"d7e1d7f0",
		16#25a4# => X"d7e1e7f4",
		16#25a5# => X"d7e1f7f8",
		16#25a6# => X"9c21fa78",
		16#25a7# => X"a9c50000",
		16#25a8# => X"d4011828",
		16#25a9# => X"d4012020",
		16#25aa# => X"04001636",
		16#25ab# => X"d401302c",
		16#25ac# => X"856b0000",
		16#25ad# => X"a86b0000",
		16#25ae# => X"07ffffaf",
		16#25af# => X"d4015848",
		16#25b0# => X"84410028",
		16#25b1# => X"bc020000",
		16#25b2# => X"10000006",
		16#25b3# => X"d4015854",
		16#25b4# => X"84420038",
		16#25b5# => X"bc220000",
		16#25b6# => X"0c00012d",
		16#25b7# => X"15000000",
		16#25b8# => X"84610020",
		16#25b9# => X"9843000c",
		16#25ba# => X"a4e2ffff",
		16#25bb# => X"a4a72000",
		16#25bc# => X"bc250000",
		16#25bd# => X"1000000b",
		16#25be# => X"a4a70008",
		16#25bf# => X"84a30064",
		16#25c0# => X"9c60dfff",
		16#25c1# => X"a8422000",
		16#25c2# => X"84810020",
		16#25c3# => X"e0a51803",
		16#25c4# => X"dc04100c",
		16#25c5# => X"d4042864",
		16#25c6# => X"a4e2ffff",
		16#25c7# => X"a4a70008",
		16#25c8# => X"bc050000",
		16#25c9# => X"1000076f",
		16#25ca# => X"84810020",
		16#25cb# => X"84a40010",
		16#25cc# => X"bc250000",
		16#25cd# => X"0c00076c",
		16#25ce# => X"84610028",
		16#25cf# => X"a4e7001a",
		16#25d0# => X"bc27000a",
		16#25d1# => X"0c0000e5",
		16#25d2# => X"84610020",
		16#25d3# => X"9c400000",
		16#25d4# => X"9c610538",
		16#25d5# => X"9c810537",
		16#25d6# => X"d4011814",
		16#25d7# => X"d4012010",
		16#25d8# => X"9c600000",
		16#25d9# => X"d4011038",
		16#25da# => X"9c4104d0",
		16#25db# => X"d4011d40",
		16#25dc# => X"d4011538",
		16#25dd# => X"d4011d3c",
		16#25de# => X"d401184c",
		16#25df# => X"d4011850",
		16#25e0# => X"d401185c",
		16#25e1# => X"d4011858",
		16#25e2# => X"d4011830",
		16#25e3# => X"aac20000",
		16#25e4# => X"84610010",
		16#25e5# => X"84410014",
		16#25e6# => X"9c810544",
		16#25e7# => X"e0421802",
		16#25e8# => X"d401701c",
		16#25e9# => X"d4011064",
		16#25ea# => X"9c41046f",
		16#25eb# => X"d4012008",
		16#25ec# => X"d401100c",
		16#25ed# => X"8461001c",
		16#25ee# => X"90a30000",
		16#25ef# => X"ac450025",
		16#25f0# => X"a44200ff",
		16#25f1# => X"bc020000",
		16#25f2# => X"100000f5",
		16#25f3# => X"a44500ff",
		16#25f4# => X"bc020000",
		16#25f5# => X"100000f2",
		16#25f6# => X"15000000",
		16#25f7# => X"00000005",
		16#25f8# => X"a9c30000",
		16#25f9# => X"bc220000",
		16#25fa# => X"0c00000a",
		16#25fb# => X"8481001c",
		16#25fc# => X"9dce0001",
		16#25fd# => X"90ae0000",
		16#25fe# => X"ac450025",
		16#25ff# => X"a44200ff",
		16#2600# => X"bc020000",
		16#2601# => X"0ffffff8",
		16#2602# => X"a44500ff",
		16#2603# => X"8481001c",
		16#2604# => X"e04e2002",
		16#2605# => X"bc020000",
		16#2606# => X"10000010",
		16#2607# => X"86410540",
		16#2608# => X"8601053c",
		16#2609# => X"e2521000",
		16#260a# => X"9e100001",
		16#260b# => X"d4162000",
		16#260c# => X"d4161004",
		16#260d# => X"d4019540",
		16#260e# => X"bd500007",
		16#260f# => X"10000080",
		16#2610# => X"d401853c",
		16#2611# => X"9ed60008",
		16#2612# => X"84610030",
		16#2613# => X"e0631000",
		16#2614# => X"d4011830",
		16#2615# => X"90ae0000",
		16#2616# => X"bc050000",
		16#2617# => X"10000081",
		16#2618# => X"9d000000",
		16#2619# => X"9dce0001",
		16#261a# => X"9c800000",
		16#261b# => X"d401701c",
		16#261c# => X"d801255b",
		16#261d# => X"9e40ffff",
		16#261e# => X"d4014034",
		16#261f# => X"d4014018",
		16#2620# => X"a8ae0000",
		16#2621# => X"93c50000",
		16#2622# => X"9ca50001",
		16#2623# => X"9c7effe0",
		16#2624# => X"bc430058",
		16#2625# => X"0c000056",
		16#2626# => X"18400001",
		16#2627# => X"d401281c",
		16#2628# => X"bc1e0000",
		16#2629# => X"1000006f",
		16#262a# => X"d801455b",
		16#262b# => X"9c800001",
		16#262c# => X"9c400000",
		16#262d# => X"9c610510",
		16#262e# => X"d4012024",
		16#262f# => X"d801f510",
		16#2630# => X"d801155b",
		16#2631# => X"ab440000",
		16#2632# => X"d4011840",
		16#2633# => X"9c400000",
		16#2634# => X"d4011044",
		16#2635# => X"84410018",
		16#2636# => X"a7820002",
		16#2637# => X"bc1c0000",
		16#2638# => X"10000006",
		16#2639# => X"84810018",
		16#263a# => X"84610024",
		16#263b# => X"9c630002",
		16#263c# => X"d4011824",
		16#263d# => X"84810018",
		16#263e# => X"a4840084",
		16#263f# => X"bc040000",
		16#2640# => X"0c00022a",
		16#2641# => X"d401203c",
		16#2642# => X"84410034",
		16#2643# => X"84610024",
		16#2644# => X"e1c21802",
		16#2645# => X"bd4e0000",
		16#2646# => X"0c000224",
		16#2647# => X"bd4e0010",
		16#2648# => X"0c0006ce",
		16#2649# => X"15000000",
		16#264a# => X"1a800001",
		16#264b# => X"d401e060",
		16#264c# => X"86410540",
		16#264d# => X"ab9a0000",
		16#264e# => X"8601053c",
		16#264f# => X"aa944060",
		16#2650# => X"9f000010",
		16#2651# => X"84410028",
		16#2652# => X"00000007",
		16#2653# => X"87410020",
		16#2654# => X"9ed60008",
		16#2655# => X"9dcefff0",
		16#2656# => X"bd4e0010",
		16#2657# => X"0c000017",
		16#2658# => X"9cf60008",
		16#2659# => X"9e100001",
		16#265a# => X"9e520010",
		16#265b# => X"d416a000",
		16#265c# => X"d416c004",
		16#265d# => X"d4019540",
		16#265e# => X"bd500007",
		16#265f# => X"0ffffff5",
		16#2660# => X"d401853c",
		16#2661# => X"a8620000",
		16#2662# => X"a89a0000",
		16#2663# => X"04001f13",
		16#2664# => X"9ca10538",
		16#2665# => X"bc2b0000",
		16#2666# => X"1000003a",
		16#2667# => X"9dcefff0",
		16#2668# => X"9ce104d8",
		16#2669# => X"9ec104d0",
		16#266a# => X"86410540",
		16#266b# => X"bd4e0010",
		16#266c# => X"13ffffed",
		16#266d# => X"8601053c",
		16#266e# => X"ab5c0000",
		16#266f# => X"87810060",
		16#2670# => X"9e100001",
		16#2671# => X"e2527000",
		16#2672# => X"d416a000",
		16#2673# => X"d4167004",
		16#2674# => X"d4019540",
		16#2675# => X"bd500007",
		16#2676# => X"10000447",
		16#2677# => X"d401853c",
		16#2678# => X"9f070008",
		16#2679# => X"000001f4",
		16#267a# => X"aac70000",
		16#267b# => X"b8630002",
		16#267c# => X"a8423eec",
		16#267d# => X"e0631000",
		16#267e# => X"84630000",
		16#267f# => X"44001800",
		16#2680# => X"15000000",
		16#2681# => X"8441002c",
		16#2682# => X"8461002c",
		16#2683# => X"84420000",
		16#2684# => X"9c630004",
		16#2685# => X"d4011034",
		16#2686# => X"bd620000",
		16#2687# => X"13ffff9a",
		16#2688# => X"d401182c",
		16#2689# => X"e0401002",
		16#268a# => X"d4011034",
		16#268b# => X"84810018",
		16#268c# => X"a8840004",
		16#268d# => X"03ffff94",
		16#268e# => X"d4012018",
		16#268f# => X"84610028",
		16#2690# => X"84810020",
		16#2691# => X"04001ee5",
		16#2692# => X"9ca10538",
		16#2693# => X"bc2b0000",
		16#2694# => X"1000000c",
		16#2695# => X"9ec104d0",
		16#2696# => X"03ffff7d",
		16#2697# => X"84610030",
		16#2698# => X"84410540",
		16#2699# => X"bc020000",
		16#269a# => X"10000007",
		16#269b# => X"84610020",
		16#269c# => X"84610028",
		16#269d# => X"84810020",
		16#269e# => X"04001ed8",
		16#269f# => X"9ca10538",
		16#26a0# => X"84610020",
		16#26a1# => X"9443000c",
		16#26a2# => X"a4420040",
		16#26a3# => X"bc020000",
		16#26a4# => X"10000005",
		16#26a5# => X"85610030",
		16#26a6# => X"9c80ffff",
		16#26a7# => X"d4012030",
		16#26a8# => X"85610030",
		16#26a9# => X"9c210588",
		16#26aa# => X"8521fffc",
		16#26ab# => X"8441ffd4",
		16#26ac# => X"85c1ffd8",
		16#26ad# => X"8601ffdc",
		16#26ae# => X"8641ffe0",
		16#26af# => X"8681ffe4",
		16#26b0# => X"86c1ffe8",
		16#26b1# => X"8701ffec",
		16#26b2# => X"8741fff0",
		16#26b3# => X"8781fff4",
		16#26b4# => X"44004800",
		16#26b5# => X"87c1fff8",
		16#26b6# => X"98e3000e",
		16#26b7# => X"bd870000",
		16#26b8# => X"13ffff1b",
		16#26b9# => X"9c80fffd",
		16#26ba# => X"9e010468",
		16#26bb# => X"e0422003",
		16#26bc# => X"85e30064",
		16#26bd# => X"85a3001c",
		16#26be# => X"85830024",
		16#26bf# => X"9d610068",
		16#26c0# => X"9d000400",
		16#26c1# => X"dc011474",
		16#26c2# => X"84610028",
		16#26c3# => X"9c400000",
		16#26c4# => X"a8900000",
		16#26c5# => X"a8ae0000",
		16#26c6# => X"84c1002c",
		16#26c7# => X"d4017ccc",
		16#26c8# => X"dc013c76",
		16#26c9# => X"d4016c84",
		16#26ca# => X"d401648c",
		16#26cb# => X"d4015c68",
		16#26cc# => X"d4015c78",
		16#26cd# => X"d4014470",
		16#26ce# => X"d401447c",
		16#26cf# => X"07fffecc",
		16#26d0# => X"d4011480",
		16#26d1# => X"e58b1000",
		16#26d2# => X"10000008",
		16#26d3# => X"d4015830",
		16#26d4# => X"84610028",
		16#26d5# => X"0400100b",
		16#26d6# => X"a8900000",
		16#26d7# => X"e42b1000",
		16#26d8# => X"100006fd",
		16#26d9# => X"9c60ffff",
		16#26da# => X"94410474",
		16#26db# => X"a4420040",
		16#26dc# => X"bc020000",
		16#26dd# => X"13ffffcb",
		16#26de# => X"84810020",
		16#26df# => X"9444000c",
		16#26e0# => X"a8420040",
		16#26e1# => X"03ffffc7",
		16#26e2# => X"dc04100c",
		16#26e3# => X"0400110b",
		16#26e4# => X"84610028",
		16#26e5# => X"03fffed4",
		16#26e6# => X"84610020",
		16#26e7# => X"85c1001c",
		16#26e8# => X"03ffff2e",
		16#26e9# => X"90ae0000",
		16#26ea# => X"84610018",
		16#26eb# => X"d401281c",
		16#26ec# => X"a8630010",
		16#26ed# => X"d801455b",
		16#26ee# => X"d4011818",
		16#26ef# => X"84810018",
		16#26f0# => X"a4e40010",
		16#26f1# => X"bc070000",
		16#26f2# => X"0c000094",
		16#26f3# => X"8441002c",
		16#26f4# => X"84610018",
		16#26f5# => X"a4e30040",
		16#26f6# => X"bc070000",
		16#26f7# => X"1000008f",
		16#26f8# => X"8441002c",
		16#26f9# => X"8481002c",
		16#26fa# => X"99c40002",
		16#26fb# => X"9c840004",
		16#26fc# => X"d401202c",
		16#26fd# => X"bd8e0000",
		16#26fe# => X"1000043e",
		16#26ff# => X"e0e07002",
		16#2700# => X"9d000001",
		16#2701# => X"e0e77004",
		16#2702# => X"b967005f",
		16#2703# => X"bd920000",
		16#2704# => X"10000005",
		16#2705# => X"84610018",
		16#2706# => X"9c80ff7f",
		16#2707# => X"e0632003",
		16#2708# => X"d4011818",
		16#2709# => X"e0e09002",
		16#270a# => X"e0e79004",
		16#270b# => X"bd870000",
		16#270c# => X"10000006",
		16#270d# => X"bc080001",
		16#270e# => X"bc0b0000",
		16#270f# => X"10000260",
		16#2710# => X"bc280000",
		16#2711# => X"bc080001",
		16#2712# => X"10000395",
		16#2713# => X"bc080002",
		16#2714# => X"10000384",
		16#2715# => X"9c410538",
		16#2716# => X"d4011040",
		16#2717# => X"a8620000",
		16#2718# => X"a44e0007",
		16#2719# => X"9c63ffff",
		16#271a# => X"9d020030",
		16#271b# => X"b9ce0043",
		16#271c# => X"bc2e0000",
		16#271d# => X"13fffffb",
		16#271e# => X"d8034000",
		16#271f# => X"d4011840",
		16#2720# => X"84610018",
		16#2721# => X"a4e30001",
		16#2722# => X"bc270000",
		16#2723# => X"10000410",
		16#2724# => X"bc280030",
		16#2725# => X"84810014",
		16#2726# => X"84410040",
		16#2727# => X"e3441002",
		16#2728# => X"e57a9000",
		16#2729# => X"10000003",
		16#272a# => X"d401d024",
		16#272b# => X"d4019024",
		16#272c# => X"9101055b",
		16#272d# => X"d4019044",
		16#272e# => X"bc080000",
		16#272f# => X"13ffff07",
		16#2730# => X"84410018",
		16#2731# => X"84810024",
		16#2732# => X"9c840001",
		16#2733# => X"03ffff02",
		16#2734# => X"d4012024",
		16#2735# => X"d801455b",
		16#2736# => X"d401281c",
		16#2737# => X"8441002c",
		16#2738# => X"8461002c",
		16#2739# => X"84420000",
		16#273a# => X"8481002c",
		16#273b# => X"d401104c",
		16#273c# => X"9c840008",
		16#273d# => X"84630004",
		16#273e# => X"8581004c",
		16#273f# => X"d4011850",
		16#2740# => X"a8ec0000",
		16#2741# => X"85610050",
		16#2742# => X"d401202c",
		16#2743# => X"a90b0000",
		16#2744# => X"e0670004",
		16#2745# => X"e0880004",
		16#2746# => X"04001d30",
		16#2747# => X"aa9e0000",
		16#2748# => X"bc2b0001",
		16#2749# => X"10000408",
		16#274a# => X"85a1004c",
		16#274b# => X"84a1004c",
		16#274c# => X"85610050",
		16#274d# => X"18400001",
		16#274e# => X"a8e50000",
		16#274f# => X"a90b0000",
		16#2750# => X"a8423ee4",
		16#2751# => X"e0670004",
		16#2752# => X"e0880004",
		16#2753# => X"84a20000",
		16#2754# => X"84c20004",
		16#2755# => X"07fff512",
		16#2756# => X"15000000",
		16#2757# => X"bd8b0000",
		16#2758# => X"10000572",
		16#2759# => X"9c60002d",
		16#275a# => X"9101055b",
		16#275b# => X"18800001",
		16#275c# => X"bd5e0047",
		16#275d# => X"a8843eaa",
		16#275e# => X"10000005",
		16#275f# => X"d4012040",
		16#2760# => X"18400001",
		16#2761# => X"a8423ea6",
		16#2762# => X"d4011040",
		16#2763# => X"9c600003",
		16#2764# => X"84810018",
		16#2765# => X"9c40ff7f",
		16#2766# => X"d4011824",
		16#2767# => X"e0841003",
		16#2768# => X"ab430000",
		16#2769# => X"9c600000",
		16#276a# => X"d4012018",
		16#276b# => X"03ffffc3",
		16#276c# => X"d4011844",
		16#276d# => X"84810018",
		16#276e# => X"a8840008",
		16#276f# => X"03fffeb2",
		16#2770# => X"d4012018",
		16#2771# => X"8441002c",
		16#2772# => X"d401281c",
		16#2773# => X"84a20000",
		16#2774# => X"9c420004",
		16#2775# => X"9c600001",
		16#2776# => X"9c800000",
		16#2777# => X"d401102c",
		16#2778# => X"9c410510",
		16#2779# => X"d4011824",
		16#277a# => X"d8012d10",
		16#277b# => X"d801255b",
		16#277c# => X"ab430000",
		16#277d# => X"03fffeb6",
		16#277e# => X"d4011040",
		16#277f# => X"84810018",
		16#2780# => X"d401281c",
		16#2781# => X"a4e40010",
		16#2782# => X"bc070000",
		16#2783# => X"13ffff71",
		16#2784# => X"d801455b",
		16#2785# => X"8441002c",
		16#2786# => X"85c20000",
		16#2787# => X"9c420004",
		16#2788# => X"03ffff75",
		16#2789# => X"d401102c",
		16#278a# => X"bc280000",
		16#278b# => X"13fffe96",
		16#278c# => X"15000000",
		16#278d# => X"03fffe94",
		16#278e# => X"9d000020",
		16#278f# => X"84810018",
		16#2790# => X"a8840001",
		16#2791# => X"03fffe90",
		16#2792# => X"d4012018",
		16#2793# => X"03fffe8e",
		16#2794# => X"9d00002b",
		16#2795# => X"84610018",
		16#2796# => X"a8630080",
		16#2797# => X"03fffe8a",
		16#2798# => X"d4011818",
		16#2799# => X"9c400000",
		16#279a# => X"9c9effd0",
		16#279b# => X"b8620003",
		16#279c# => X"e0421000",
		16#279d# => X"93c50000",
		16#279e# => X"e0421800",
		16#279f# => X"e0441000",
		16#27a0# => X"9c9effd0",
		16#27a1# => X"bca40009",
		16#27a2# => X"13fffff9",
		16#27a3# => X"9ca50001",
		16#27a4# => X"03fffe7f",
		16#27a5# => X"d4011034",
		16#27a6# => X"93c50000",
		16#27a7# => X"bc1e002a",
		16#27a8# => X"1000061d",
		16#27a9# => X"9ca50001",
		16#27aa# => X"9c9effd0",
		16#27ab# => X"bca40009",
		16#27ac# => X"0c00000b",
		16#27ad# => X"9e400000",
		16#27ae# => X"b8520003",
		16#27af# => X"e2529000",
		16#27b0# => X"93c50000",
		16#27b1# => X"e2521000",
		16#27b2# => X"e2522000",
		16#27b3# => X"9c9effd0",
		16#27b4# => X"bca40009",
		16#27b5# => X"13fffff9",
		16#27b6# => X"9ca50001",
		16#27b7# => X"bd720000",
		16#27b8# => X"13fffe6c",
		16#27b9# => X"9c7effe0",
		16#27ba# => X"03fffe6a",
		16#27bb# => X"9e40ffff",
		16#27bc# => X"84410018",
		16#27bd# => X"a8420040",
		16#27be# => X"03fffe63",
		16#27bf# => X"d4011018",
		16#27c0# => X"84610018",
		16#27c1# => X"a8630010",
		16#27c2# => X"03fffe5f",
		16#27c3# => X"d4011818",
		16#27c4# => X"84410018",
		16#27c5# => X"d401281c",
		16#27c6# => X"a4a20010",
		16#27c7# => X"bc050000",
		16#27c8# => X"10000451",
		16#27c9# => X"d801455b",
		16#27ca# => X"8461002c",
		16#27cb# => X"84810030",
		16#27cc# => X"84430000",
		16#27cd# => X"9c630004",
		16#27ce# => X"d401182c",
		16#27cf# => X"03fffe1e",
		16#27d0# => X"d4022000",
		16#27d1# => X"8481002c",
		16#27d2# => X"84410018",
		16#27d3# => X"85c40000",
		16#27d4# => X"a8420002",
		16#27d5# => X"9c600030",
		16#27d6# => X"e0e07002",
		16#27d7# => X"d4011018",
		16#27d8# => X"d8011d58",
		16#27d9# => X"8441002c",
		16#27da# => X"18600001",
		16#27db# => X"e0e77004",
		16#27dc# => X"9c800078",
		16#27dd# => X"9c420004",
		16#27de# => X"a8633ec7",
		16#27df# => X"b967005f",
		16#27e0# => X"d401281c",
		16#27e1# => X"d8012559",
		16#27e2# => X"d401102c",
		16#27e3# => X"d401185c",
		16#27e4# => X"9d000002",
		16#27e5# => X"9fc00078",
		16#27e6# => X"9c400000",
		16#27e7# => X"03ffff1c",
		16#27e8# => X"d801155b",
		16#27e9# => X"9c800000",
		16#27ea# => X"8441002c",
		16#27eb# => X"d801255b",
		16#27ec# => X"d401281c",
		16#27ed# => X"84620000",
		16#27ee# => X"9dc20004",
		16#27ef# => X"bc230000",
		16#27f0# => X"0c00053b",
		16#27f1# => X"d4011840",
		16#27f2# => X"bd920000",
		16#27f3# => X"10000518",
		16#27f4# => X"84610040",
		16#27f5# => X"9c800000",
		16#27f6# => X"04001475",
		16#27f7# => X"a8b20000",
		16#27f8# => X"bc2b0000",
		16#27f9# => X"0c000597",
		16#27fa# => X"84410040",
		16#27fb# => X"e34b1002",
		16#27fc# => X"e5ba9000",
		16#27fd# => X"100004ad",
		16#27fe# => X"ac5affff",
		16#27ff# => X"9c600000",
		16#2800# => X"d4019024",
		16#2801# => X"9101055b",
		16#2802# => X"ab520000",
		16#2803# => X"d401702c",
		16#2804# => X"03ffff2a",
		16#2805# => X"d4011844",
		16#2806# => X"18600001",
		16#2807# => X"84810018",
		16#2808# => X"a8633ec7",
		16#2809# => X"a4e40010",
		16#280a# => X"d401281c",
		16#280b# => X"d801455b",
		16#280c# => X"bc070000",
		16#280d# => X"0c00003c",
		16#280e# => X"d401185c",
		16#280f# => X"84610018",
		16#2810# => X"a4e30040",
		16#2811# => X"bc070000",
		16#2812# => X"10000038",
		16#2813# => X"8441002c",
		16#2814# => X"8481002c",
		16#2815# => X"85c40000",
		16#2816# => X"9c840004",
		16#2817# => X"a5ceffff",
		16#2818# => X"e0e07002",
		16#2819# => X"e0e77004",
		16#281a# => X"b967005f",
		16#281b# => X"bc0b0000",
		16#281c# => X"10000036",
		16#281d# => X"d401202c",
		16#281e# => X"84610018",
		16#281f# => X"a5030001",
		16#2820# => X"bc080000",
		16#2821# => X"10000031",
		16#2822# => X"9c800030",
		16#2823# => X"a8630002",
		16#2824# => X"d8012558",
		16#2825# => X"d801f559",
		16#2826# => X"d4011818",
		16#2827# => X"9d600001",
		16#2828# => X"03ffffbe",
		16#2829# => X"9d000002",
		16#282a# => X"84810018",
		16#282b# => X"a8840010",
		16#282c# => X"03fffdf5",
		16#282d# => X"d4012018",
		16#282e# => X"84610018",
		16#282f# => X"d401281c",
		16#2830# => X"a8630010",
		16#2831# => X"d4011818",
		16#2832# => X"84810018",
		16#2833# => X"a4e40010",
		16#2834# => X"bc070000",
		16#2835# => X"100002b7",
		16#2836# => X"84610018",
		16#2837# => X"8441002c",
		16#2838# => X"9d000001",
		16#2839# => X"85c20000",
		16#283a# => X"9c420004",
		16#283b# => X"e0e07002",
		16#283c# => X"d401102c",
		16#283d# => X"e0e77004",
		16#283e# => X"03ffffa8",
		16#283f# => X"b967005f",
		16#2840# => X"18600001",
		16#2841# => X"84810018",
		16#2842# => X"a8633eb6",
		16#2843# => X"a4e40010",
		16#2844# => X"d401281c",
		16#2845# => X"d801455b",
		16#2846# => X"bc070000",
		16#2847# => X"13ffffc8",
		16#2848# => X"d401185c",
		16#2849# => X"8441002c",
		16#284a# => X"85c20000",
		16#284b# => X"9c420004",
		16#284c# => X"e0e07002",
		16#284d# => X"e0e77004",
		16#284e# => X"b967005f",
		16#284f# => X"bc0b0000",
		16#2850# => X"0fffffce",
		16#2851# => X"d401102c",
		16#2852# => X"03ffff94",
		16#2853# => X"9d000002",
		16#2854# => X"84810018",
		16#2855# => X"d401281c",
		16#2856# => X"a8840010",
		16#2857# => X"d4012018",
		16#2858# => X"84410018",
		16#2859# => X"a5020010",
		16#285a# => X"bc080000",
		16#285b# => X"1000029e",
		16#285c# => X"84810018",
		16#285d# => X"8461002c",
		16#285e# => X"9d000000",
		16#285f# => X"85c30000",
		16#2860# => X"9c630004",
		16#2861# => X"e0e07002",
		16#2862# => X"d401182c",
		16#2863# => X"e0e77004",
		16#2864# => X"03ffff82",
		16#2865# => X"b967005f",
		16#2866# => X"03fffff2",
		16#2867# => X"d401281c",
		16#2868# => X"03ffffca",
		16#2869# => X"d401281c",
		16#286a# => X"9f160008",
		16#286b# => X"86410540",
		16#286c# => X"8601053c",
		16#286d# => X"9041055b",
		16#286e# => X"bc020000",
		16#286f# => X"1000000f",
		16#2870# => X"bc1c0000",
		16#2871# => X"9e100001",
		16#2872# => X"9e520001",
		16#2873# => X"9c81055b",
		16#2874# => X"9c400001",
		16#2875# => X"d4162000",
		16#2876# => X"d4161004",
		16#2877# => X"d4019540",
		16#2878# => X"bd500007",
		16#2879# => X"100001d0",
		16#287a# => X"d401853c",
		16#287b# => X"aad80000",
		16#287c# => X"9f180008",
		16#287d# => X"bc1c0000",
		16#287e# => X"1000000f",
		16#287f# => X"8441003c",
		16#2880# => X"9e100001",
		16#2881# => X"9e520002",
		16#2882# => X"9c610558",
		16#2883# => X"9c800002",
		16#2884# => X"d4161800",
		16#2885# => X"d4162004",
		16#2886# => X"d4019540",
		16#2887# => X"bd500007",
		16#2888# => X"100001cc",
		16#2889# => X"d401853c",
		16#288a# => X"aad80000",
		16#288b# => X"9f180008",
		16#288c# => X"8441003c",
		16#288d# => X"bc220080",
		16#288e# => X"0c0000ee",
		16#288f# => X"84610034",
		16#2890# => X"84610044",
		16#2891# => X"e043d002",
		16#2892# => X"bda20000",
		16#2893# => X"1000002e",
		16#2894# => X"bda20010",
		16#2895# => X"100003c5",
		16#2896# => X"15000000",
		16#2897# => X"1a800001",
		16#2898# => X"9dc00010",
		16#2899# => X"aa944050",
		16#289a# => X"87010028",
		16#289b# => X"00000007",
		16#289c# => X"87810020",
		16#289d# => X"9ed60008",
		16#289e# => X"9c42fff0",
		16#289f# => X"bd420010",
		16#28a0# => X"0c000017",
		16#28a1# => X"9cb60008",
		16#28a2# => X"9e100001",
		16#28a3# => X"9e520010",
		16#28a4# => X"d416a000",
		16#28a5# => X"d4167004",
		16#28a6# => X"d4019540",
		16#28a7# => X"bd500007",
		16#28a8# => X"0ffffff5",
		16#28a9# => X"d401853c",
		16#28aa# => X"a8780000",
		16#28ab# => X"a89c0000",
		16#28ac# => X"04001cca",
		16#28ad# => X"9ca10538",
		16#28ae# => X"bc2b0000",
		16#28af# => X"13fffdf1",
		16#28b0# => X"9c42fff0",
		16#28b1# => X"9ca104d8",
		16#28b2# => X"9ec104d0",
		16#28b3# => X"86410540",
		16#28b4# => X"bd420010",
		16#28b5# => X"13ffffed",
		16#28b6# => X"8601053c",
		16#28b7# => X"9e100001",
		16#28b8# => X"e2521000",
		16#28b9# => X"d416a000",
		16#28ba# => X"d4161004",
		16#28bb# => X"d4019540",
		16#28bc# => X"bd500007",
		16#28bd# => X"10000181",
		16#28be# => X"d401853c",
		16#28bf# => X"9f050008",
		16#28c0# => X"aac50000",
		16#28c1# => X"84810018",
		16#28c2# => X"a4440100",
		16#28c3# => X"bc220000",
		16#28c4# => X"10000054",
		16#28c5# => X"bdbe0065",
		16#28c6# => X"9e100001",
		16#28c7# => X"e252d000",
		16#28c8# => X"84410040",
		16#28c9# => X"d416d004",
		16#28ca# => X"d4161000",
		16#28cb# => X"d4019540",
		16#28cc# => X"bdb00007",
		16#28cd# => X"0c00010c",
		16#28ce# => X"d401853c",
		16#28cf# => X"84810018",
		16#28d0# => X"a4440004",
		16#28d1# => X"bc220000",
		16#28d2# => X"0c000039",
		16#28d3# => X"84410024",
		16#28d4# => X"84410034",
		16#28d5# => X"84610024",
		16#28d6# => X"e1c21802",
		16#28d7# => X"bd4e0000",
		16#28d8# => X"0c000032",
		16#28d9# => X"bdae0010",
		16#28da# => X"10000468",
		16#28db# => X"15000000",
		16#28dc# => X"1a800001",
		16#28dd# => X"8601053c",
		16#28de# => X"aa944060",
		16#28df# => X"9ec00010",
		16#28e0# => X"84410028",
		16#28e1# => X"00000006",
		16#28e2# => X"87410020",
		16#28e3# => X"9dcefff0",
		16#28e4# => X"bd4e0010",
		16#28e5# => X"0c000016",
		16#28e6# => X"9f180008",
		16#28e7# => X"9e100001",
		16#28e8# => X"9e520010",
		16#28e9# => X"d418a000",
		16#28ea# => X"d418b004",
		16#28eb# => X"d4019540",
		16#28ec# => X"bd500007",
		16#28ed# => X"0ffffff6",
		16#28ee# => X"d401853c",
		16#28ef# => X"a8620000",
		16#28f0# => X"a89a0000",
		16#28f1# => X"04001c85",
		16#28f2# => X"9ca10538",
		16#28f3# => X"bc2b0000",
		16#28f4# => X"13fffdac",
		16#28f5# => X"9dcefff0",
		16#28f6# => X"9f0104d0",
		16#28f7# => X"86410540",
		16#28f8# => X"bd4e0010",
		16#28f9# => X"13ffffee",
		16#28fa# => X"8601053c",
		16#28fb# => X"9e100001",
		16#28fc# => X"e24e9000",
		16#28fd# => X"d418a000",
		16#28fe# => X"d4187004",
		16#28ff# => X"d4019540",
		16#2900# => X"bdb00007",
		16#2901# => X"10000009",
		16#2902# => X"d401853c",
		16#2903# => X"84610028",
		16#2904# => X"84810020",
		16#2905# => X"04001c71",
		16#2906# => X"9ca10538",
		16#2907# => X"bc2b0000",
		16#2908# => X"13fffd98",
		16#2909# => X"86410540",
		16#290a# => X"84410024",
		16#290b# => X"84810034",
		16#290c# => X"e5622000",
		16#290d# => X"10000003",
		16#290e# => X"84610030",
		16#290f# => X"a8440000",
		16#2910# => X"bc120000",
		16#2911# => X"e0631000",
		16#2912# => X"0c00009c",
		16#2913# => X"d4011830",
		16#2914# => X"9c800000",
		16#2915# => X"9ec104d0",
		16#2916# => X"03fffcd7",
		16#2917# => X"d401253c",
		16#2918# => X"100000ca",
		16#2919# => X"84410038",
		16#291a# => X"84a1004c",
		16#291b# => X"85810050",
		16#291c# => X"18600001",
		16#291d# => X"a8e50000",
		16#291e# => X"a8633ee4",
		16#291f# => X"a90c0000",
		16#2920# => X"84a30000",
		16#2921# => X"84c30004",
		16#2922# => X"e0670004",
		16#2923# => X"e0880004",
		16#2924# => X"07fff2cb",
		16#2925# => X"15000000",
		16#2926# => X"bc0b0000",
		16#2927# => X"0c000138",
		16#2928# => X"85c10554",
		16#2929# => X"18a00001",
		16#292a# => X"9e100001",
		16#292b# => X"9e520001",
		16#292c# => X"a8a53edf",
		16#292d# => X"9c800001",
		16#292e# => X"d4162800",
		16#292f# => X"d4162004",
		16#2930# => X"d4019540",
		16#2931# => X"bdb00007",
		16#2932# => X"0c00032c",
		16#2933# => X"d401853c",
		16#2934# => X"84a10554",
		16#2935# => X"84410038",
		16#2936# => X"e5851000",
		16#2937# => X"10000006",
		16#2938# => X"84610018",
		16#2939# => X"a4a30001",
		16#293a# => X"bc050000",
		16#293b# => X"13ffff95",
		16#293c# => X"84810018",
		16#293d# => X"8601053c",
		16#293e# => X"84810054",
		16#293f# => X"9e100001",
		16#2940# => X"e2522000",
		16#2941# => X"84410048",
		16#2942# => X"d4182004",
		16#2943# => X"d4181000",
		16#2944# => X"d4019540",
		16#2945# => X"bd500007",
		16#2946# => X"100003ac",
		16#2947# => X"d401853c",
		16#2948# => X"9cb80008",
		16#2949# => X"84610038",
		16#294a# => X"9dc3ffff",
		16#294b# => X"bdae0000",
		16#294c# => X"100003af",
		16#294d# => X"bd4e0010",
		16#294e# => X"0c0001f6",
		16#294f# => X"1a800001",
		16#2950# => X"8601053c",
		16#2951# => X"aa944050",
		16#2952# => X"9ec00010",
		16#2953# => X"84410028",
		16#2954# => X"00000008",
		16#2955# => X"87410020",
		16#2956# => X"9ca50008",
		16#2957# => X"9f050008",
		16#2958# => X"9dcefff0",
		16#2959# => X"bd4e0010",
		16#295a# => X"0c0001ed",
		16#295b# => X"15000000",
		16#295c# => X"9e100001",
		16#295d# => X"9e520010",
		16#295e# => X"d405a000",
		16#295f# => X"d405b004",
		16#2960# => X"d4019540",
		16#2961# => X"bd500007",
		16#2962# => X"0ffffff4",
		16#2963# => X"d401853c",
		16#2964# => X"a8620000",
		16#2965# => X"a89a0000",
		16#2966# => X"04001c10",
		16#2967# => X"9ca10538",
		16#2968# => X"bc2b0000",
		16#2969# => X"13fffd37",
		16#296a# => X"9f0104d8",
		16#296b# => X"9ca104d0",
		16#296c# => X"86410540",
		16#296d# => X"03ffffeb",
		16#296e# => X"8601053c",
		16#296f# => X"100000cc",
		16#2970# => X"9c410538",
		16#2971# => X"84410018",
		16#2972# => X"a4e20001",
		16#2973# => X"bc070000",
		16#2974# => X"10000121",
		16#2975# => X"9c610538",
		16#2976# => X"9c600030",
		16#2977# => X"9c810537",
		16#2978# => X"d8011d37",
		16#2979# => X"87410064",
		16#297a# => X"03fffdae",
		16#297b# => X"d4012040",
		16#297c# => X"84810024",
		16#297d# => X"e1c32002",
		16#297e# => X"bd4e0000",
		16#297f# => X"0c000186",
		16#2980# => X"bdae0010",
		16#2981# => X"1000040b",
		16#2982# => X"15000000",
		16#2983# => X"1a800001",
		16#2984# => X"9f000010",
		16#2985# => X"aa944050",
		16#2986# => X"84410028",
		16#2987# => X"00000007",
		16#2988# => X"87810020",
		16#2989# => X"9ed60008",
		16#298a# => X"9dcefff0",
		16#298b# => X"bd4e0010",
		16#298c# => X"0c000017",
		16#298d# => X"9d160008",
		16#298e# => X"9e100001",
		16#298f# => X"9e520010",
		16#2990# => X"d416a000",
		16#2991# => X"d416c004",
		16#2992# => X"d4019540",
		16#2993# => X"bd500007",
		16#2994# => X"0ffffff5",
		16#2995# => X"d401853c",
		16#2996# => X"a8620000",
		16#2997# => X"a89c0000",
		16#2998# => X"04001bde",
		16#2999# => X"9ca10538",
		16#299a# => X"bc2b0000",
		16#299b# => X"13fffd05",
		16#299c# => X"9dcefff0",
		16#299d# => X"9d0104d8",
		16#299e# => X"9ec104d0",
		16#299f# => X"86410540",
		16#29a0# => X"bd4e0010",
		16#29a1# => X"13ffffed",
		16#29a2# => X"8601053c",
		16#29a3# => X"9e100001",
		16#29a4# => X"e2527000",
		16#29a5# => X"d416a000",
		16#29a6# => X"d4167004",
		16#29a7# => X"d4019540",
		16#29a8# => X"bd500007",
		16#29a9# => X"1000017f",
		16#29aa# => X"d401853c",
		16#29ab# => X"9f080008",
		16#29ac# => X"03fffee4",
		16#29ad# => X"aac80000",
		16#29ae# => X"84610028",
		16#29af# => X"84810020",
		16#29b0# => X"04001bc6",
		16#29b1# => X"9ca10538",
		16#29b2# => X"bc2b0000",
		16#29b3# => X"0fffff62",
		16#29b4# => X"9c800000",
		16#29b5# => X"03fffcec",
		16#29b6# => X"84610020",
		16#29b7# => X"9e100001",
		16#29b8# => X"84410040",
		16#29b9# => X"d4161000",
		16#29ba# => X"d4167004",
		16#29bb# => X"d4015d40",
		16#29bc# => X"d401853c",
		16#29bd# => X"bdb00007",
		16#29be# => X"0c000388",
		16#29bf# => X"a84e0000",
		16#29c0# => X"84610054",
		16#29c1# => X"9e100001",
		16#29c2# => X"e16b1800",
		16#29c3# => X"84810048",
		16#29c4# => X"d4181804",
		16#29c5# => X"d4182000",
		16#29c6# => X"d4015d40",
		16#29c7# => X"bd500007",
		16#29c8# => X"10000391",
		16#29c9# => X"d401853c",
		16#29ca# => X"9f180008",
		16#29cb# => X"84610038",
		16#29cc# => X"86410540",
		16#29cd# => X"e1c37002",
		16#29ce# => X"8601053c",
		16#29cf# => X"84810040",
		16#29d0# => X"9e100001",
		16#29d1# => X"e1041000",
		16#29d2# => X"e2527000",
		16#29d3# => X"d4184000",
		16#29d4# => X"d4187004",
		16#29d5# => X"d4019540",
		16#29d6# => X"bd500007",
		16#29d7# => X"0c000281",
		16#29d8# => X"d401853c",
		16#29d9# => X"84610028",
		16#29da# => X"84810020",
		16#29db# => X"04001b9b",
		16#29dc# => X"9ca10538",
		16#29dd# => X"bc2b0000",
		16#29de# => X"13fffcc2",
		16#29df# => X"9f0104d0",
		16#29e0# => X"03fffeef",
		16#29e1# => X"86410540",
		16#29e2# => X"bd420001",
		16#29e3# => X"0c000040",
		16#29e4# => X"84610018",
		16#29e5# => X"9e100001",
		16#29e6# => X"9e520001",
		16#29e7# => X"84810040",
		16#29e8# => X"9c400001",
		16#29e9# => X"d4162000",
		16#29ea# => X"d4161004",
		16#29eb# => X"d4019540",
		16#29ec# => X"bd500007",
		16#29ed# => X"1000011a",
		16#29ee# => X"d401853c",
		16#29ef# => X"9dd80008",
		16#29f0# => X"84610054",
		16#29f1# => X"9e100001",
		16#29f2# => X"e2521800",
		16#29f3# => X"84810048",
		16#29f4# => X"d4181804",
		16#29f5# => X"d4182000",
		16#29f6# => X"d4019540",
		16#29f7# => X"bd500007",
		16#29f8# => X"1000011a",
		16#29f9# => X"d401853c",
		16#29fa# => X"9f4e0008",
		16#29fb# => X"84a1004c",
		16#29fc# => X"85810050",
		16#29fd# => X"18400001",
		16#29fe# => X"a8e50000",
		16#29ff# => X"a90c0000",
		16#2a00# => X"a8423ee4",
		16#2a01# => X"e0670004",
		16#2a02# => X"e0880004",
		16#2a03# => X"84a20000",
		16#2a04# => X"84c20004",
		16#2a05# => X"07fff208",
		16#2a06# => X"15000000",
		16#2a07# => X"bc2b0000",
		16#2a08# => X"0c0000c0",
		16#2a09# => X"84410038",
		16#2a0a# => X"84610038",
		16#2a0b# => X"84810040",
		16#2a0c# => X"9d03ffff",
		16#2a0d# => X"9e100001",
		16#2a0e# => X"9ca40001",
		16#2a0f# => X"e2524000",
		16#2a10# => X"d40e2800",
		16#2a11# => X"d40e4004",
		16#2a12# => X"d4019540",
		16#2a13# => X"bd500007",
		16#2a14# => X"1000001c",
		16#2a15# => X"d401853c",
		16#2a16# => X"9f1a0008",
		16#2a17# => X"84410058",
		16#2a18# => X"9e100001",
		16#2a19# => X"e2521000",
		16#2a1a# => X"9c610544",
		16#2a1b# => X"d41a1004",
		16#2a1c# => X"d41a1800",
		16#2a1d# => X"d4019540",
		16#2a1e# => X"bdb00007",
		16#2a1f# => X"13fffeb0",
		16#2a20# => X"d401853c",
		16#2a21# => X"03ffffb9",
		16#2a22# => X"84610028",
		16#2a23# => X"a4a30001",
		16#2a24# => X"bc050000",
		16#2a25# => X"0fffffc0",
		16#2a26# => X"84610040",
		16#2a27# => X"9e100001",
		16#2a28# => X"9e520001",
		16#2a29# => X"9c800001",
		16#2a2a# => X"d4161800",
		16#2a2b# => X"d4162004",
		16#2a2c# => X"d4019540",
		16#2a2d# => X"bd500007",
		16#2a2e# => X"0c00029f",
		16#2a2f# => X"d401853c",
		16#2a30# => X"84610028",
		16#2a31# => X"84810020",
		16#2a32# => X"04001b44",
		16#2a33# => X"9ca10538",
		16#2a34# => X"bc2b0000",
		16#2a35# => X"13fffc6b",
		16#2a36# => X"9f0104d8",
		16#2a37# => X"9f4104d0",
		16#2a38# => X"86410540",
		16#2a39# => X"03ffffde",
		16#2a3a# => X"8601053c",
		16#2a3b# => X"ab4b0000",
		16#2a3c# => X"03fffcec",
		16#2a3d# => X"d4011040",
		16#2a3e# => X"84610028",
		16#2a3f# => X"84810020",
		16#2a40# => X"04001b36",
		16#2a41# => X"9ca10538",
		16#2a42# => X"bc2b0000",
		16#2a43# => X"13fffc5d",
		16#2a44# => X"9f0104d8",
		16#2a45# => X"9ec104d0",
		16#2a46# => X"86410540",
		16#2a47# => X"03fffe7a",
		16#2a48# => X"8601053c",
		16#2a49# => X"84610028",
		16#2a4a# => X"84810020",
		16#2a4b# => X"04001b2b",
		16#2a4c# => X"9ca10538",
		16#2a4d# => X"bc2b0000",
		16#2a4e# => X"13fffc52",
		16#2a4f# => X"9f0104d8",
		16#2a50# => X"9ec104d0",
		16#2a51# => X"86410540",
		16#2a52# => X"03fffe2b",
		16#2a53# => X"8601053c",
		16#2a54# => X"84610028",
		16#2a55# => X"84810020",
		16#2a56# => X"04001b20",
		16#2a57# => X"9ca10538",
		16#2a58# => X"bc2b0000",
		16#2a59# => X"13fffc47",
		16#2a5a# => X"9f0104d8",
		16#2a5b# => X"9ec104d0",
		16#2a5c# => X"86410540",
		16#2a5d# => X"03fffe2f",
		16#2a5e# => X"8601053c",
		16#2a5f# => X"bd4e0000",
		16#2a60# => X"0c000207",
		16#2a61# => X"84410038",
		16#2a62# => X"e58e1000",
		16#2a63# => X"13ffff54",
		16#2a64# => X"e16e9000",
		16#2a65# => X"9e100001",
		16#2a66# => X"e2521000",
		16#2a67# => X"84610040",
		16#2a68# => X"d4161004",
		16#2a69# => X"d4161800",
		16#2a6a# => X"d4019540",
		16#2a6b# => X"bdb00007",
		16#2a6c# => X"0c0002f6",
		16#2a6d# => X"d401853c",
		16#2a6e# => X"84810038",
		16#2a6f# => X"e1ce2002",
		16#2a70# => X"bdae0000",
		16#2a71# => X"100001d7",
		16#2a72# => X"bd4e0010",
		16#2a73# => X"0c0001c1",
		16#2a74# => X"1a800001",
		16#2a75# => X"a8b80000",
		16#2a76# => X"8601053c",
		16#2a77# => X"aa944050",
		16#2a78# => X"9ec00010",
		16#2a79# => X"84410028",
		16#2a7a# => X"00000008",
		16#2a7b# => X"87410020",
		16#2a7c# => X"9ca50008",
		16#2a7d# => X"9f050008",
		16#2a7e# => X"9dcefff0",
		16#2a7f# => X"bd4e0010",
		16#2a80# => X"0c0001b8",
		16#2a81# => X"15000000",
		16#2a82# => X"9e100001",
		16#2a83# => X"9e520010",
		16#2a84# => X"d405a000",
		16#2a85# => X"d405b004",
		16#2a86# => X"d4019540",
		16#2a87# => X"bd500007",
		16#2a88# => X"0ffffff4",
		16#2a89# => X"d401853c",
		16#2a8a# => X"a8620000",
		16#2a8b# => X"a89a0000",
		16#2a8c# => X"04001aea",
		16#2a8d# => X"9ca10538",
		16#2a8e# => X"bc2b0000",
		16#2a8f# => X"13fffc11",
		16#2a90# => X"9f0104d8",
		16#2a91# => X"9ca104d0",
		16#2a92# => X"86410540",
		16#2a93# => X"03ffffeb",
		16#2a94# => X"8601053c",
		16#2a95# => X"ab480000",
		16#2a96# => X"03fffc92",
		16#2a97# => X"d4011840",
		16#2a98# => X"9c610538",
		16#2a99# => X"8481005c",
		16#2a9a# => X"d4011840",
		16#2a9b# => X"a44e000f",
		16#2a9c# => X"9c63ffff",
		16#2a9d# => X"e0441000",
		16#2a9e# => X"b9ce0044",
		16#2a9f# => X"8c420000",
		16#2aa0# => X"bc2e0000",
		16#2aa1# => X"13fffffa",
		16#2aa2# => X"d8031000",
		16#2aa3# => X"84810014",
		16#2aa4# => X"d4011840",
		16#2aa5# => X"03fffc83",
		16#2aa6# => X"e3441802",
		16#2aa7# => X"bc4e0009",
		16#2aa8# => X"0c00000e",
		16#2aa9# => X"9e010538",
		16#2aaa# => X"a86e0000",
		16#2aab# => X"9c80000a",
		16#2aac# => X"0400239a",
		16#2aad# => X"9e10ffff",
		16#2aae# => X"9d6b0030",
		16#2aaf# => X"a86e0000",
		16#2ab0# => X"9c80000a",
		16#2ab1# => X"07ffe810",
		16#2ab2# => X"d8105800",
		16#2ab3# => X"bc4b0009",
		16#2ab4# => X"13fffff6",
		16#2ab5# => X"a9cb0000",
		16#2ab6# => X"9e10ffff",
		16#2ab7# => X"84410014",
		16#2ab8# => X"9dce0030",
		16#2ab9# => X"d4018040",
		16#2aba# => X"e3428002",
		16#2abb# => X"03fffc6d",
		16#2abc# => X"d8107000",
		16#2abd# => X"84610028",
		16#2abe# => X"84810020",
		16#2abf# => X"04001ab7",
		16#2ac0# => X"9ca10538",
		16#2ac1# => X"bc2b0000",
		16#2ac2# => X"13fffbde",
		16#2ac3# => X"9f0104d8",
		16#2ac4# => X"9ec104d0",
		16#2ac5# => X"86410540",
		16#2ac6# => X"03fffda7",
		16#2ac7# => X"8601053c",
		16#2ac8# => X"9ec2ffff",
		16#2ac9# => X"bd560000",
		16#2aca# => X"0c000225",
		16#2acb# => X"bdb60010",
		16#2acc# => X"10000051",
		16#2acd# => X"1a800001",
		16#2ace# => X"9f000010",
		16#2acf# => X"aa944050",
		16#2ad0# => X"84410028",
		16#2ad1# => X"00000008",
		16#2ad2# => X"87810020",
		16#2ad3# => X"9dce0008",
		16#2ad4# => X"9f4e0008",
		16#2ad5# => X"9ed6fff0",
		16#2ad6# => X"bd560010",
		16#2ad7# => X"0c000047",
		16#2ad8# => X"15000000",
		16#2ad9# => X"9e100001",
		16#2ada# => X"9e520010",
		16#2adb# => X"d40ea000",
		16#2adc# => X"d40ec004",
		16#2add# => X"d4019540",
		16#2ade# => X"bd500007",
		16#2adf# => X"0ffffff4",
		16#2ae0# => X"d401853c",
		16#2ae1# => X"a8620000",
		16#2ae2# => X"a89c0000",
		16#2ae3# => X"04001a93",
		16#2ae4# => X"9ca10538",
		16#2ae5# => X"bc2b0000",
		16#2ae6# => X"13fffbba",
		16#2ae7# => X"9f4104d8",
		16#2ae8# => X"9dc104d0",
		16#2ae9# => X"86410540",
		16#2aea# => X"03ffffeb",
		16#2aeb# => X"8601053c",
		16#2aec# => X"a4e30040",
		16#2aed# => X"bc070000",
		16#2aee# => X"10000136",
		16#2aef# => X"8441002c",
		16#2af0# => X"8481002c",
		16#2af1# => X"9d000001",
		16#2af2# => X"85c40000",
		16#2af3# => X"9c840004",
		16#2af4# => X"a5ceffff",
		16#2af5# => X"d401202c",
		16#2af6# => X"e0e07002",
		16#2af7# => X"03fffcef",
		16#2af8# => X"b967005f",
		16#2af9# => X"a5640040",
		16#2afa# => X"bc0b0000",
		16#2afb# => X"10000131",
		16#2afc# => X"8461002c",
		16#2afd# => X"8441002c",
		16#2afe# => X"85c20000",
		16#2aff# => X"9c420004",
		16#2b00# => X"a5ceffff",
		16#2b01# => X"d401102c",
		16#2b02# => X"e0e07002",
		16#2b03# => X"03fffce3",
		16#2b04# => X"b967005f",
		16#2b05# => X"03fffd8b",
		16#2b06# => X"9f160008",
		16#2b07# => X"84610028",
		16#2b08# => X"84810020",
		16#2b09# => X"04001a6d",
		16#2b0a# => X"9ca10538",
		16#2b0b# => X"bc2b0000",
		16#2b0c# => X"13fffb94",
		16#2b0d# => X"9dc104d8",
		16#2b0e# => X"9f0104d0",
		16#2b0f# => X"86410540",
		16#2b10# => X"03fffee0",
		16#2b11# => X"8601053c",
		16#2b12# => X"84610028",
		16#2b13# => X"84810020",
		16#2b14# => X"04001a62",
		16#2b15# => X"9ca10538",
		16#2b16# => X"bc2b0000",
		16#2b17# => X"13fffb89",
		16#2b18# => X"9f4104d8",
		16#2b19# => X"9dc104d0",
		16#2b1a# => X"86410540",
		16#2b1b# => X"03fffee0",
		16#2b1c# => X"8601053c",
		16#2b1d# => X"aa944050",
		16#2b1e# => X"9e100001",
		16#2b1f# => X"e252b000",
		16#2b20# => X"d40ea000",
		16#2b21# => X"d40eb004",
		16#2b22# => X"d4019540",
		16#2b23# => X"bd500007",
		16#2b24# => X"0ffffef2",
		16#2b25# => X"d401853c",
		16#2b26# => X"03ffff0b",
		16#2b27# => X"84610028",
		16#2b28# => X"84610028",
		16#2b29# => X"84810020",
		16#2b2a# => X"04001a4c",
		16#2b2b# => X"9ca10538",
		16#2b2c# => X"bc2b0000",
		16#2b2d# => X"13fffb73",
		16#2b2e# => X"9f0104d8",
		16#2b2f# => X"9ec104d0",
		16#2b30# => X"86410540",
		16#2b31# => X"03fffd5f",
		16#2b32# => X"8601053c",
		16#2b33# => X"0c0001e9",
		16#2b34# => X"84410040",
		16#2b35# => X"9c600030",
		16#2b36# => X"9c42ffff",
		16#2b37# => X"d4011040",
		16#2b38# => X"d8021800",
		16#2b39# => X"84810014",
		16#2b3a# => X"03fffbee",
		16#2b3b# => X"e3441002",
		16#2b3c# => X"e1c07002",
		16#2b3d# => X"9c60002d",
		16#2b3e# => X"e1607002",
		16#2b3f# => X"d8011d5b",
		16#2b40# => X"e0eb7004",
		16#2b41# => X"9d000001",
		16#2b42# => X"03fffbc1",
		16#2b43# => X"b967005f",
		16#2b44# => X"9f050008",
		16#2b45# => X"8601053c",
		16#2b46# => X"aa944050",
		16#2b47# => X"9e100001",
		16#2b48# => X"e2527000",
		16#2b49# => X"d405a000",
		16#2b4a# => X"d4057004",
		16#2b4b# => X"d4019540",
		16#2b4c# => X"bdb00007",
		16#2b4d# => X"13fffd82",
		16#2b4e# => X"d401853c",
		16#2b4f# => X"03fffe8b",
		16#2b50# => X"84610028",
		16#2b51# => X"85610050",
		16#2b52# => X"a8ed0000",
		16#2b53# => X"a90b0000",
		16#2b54# => X"e0670004",
		16#2b55# => X"e0880004",
		16#2b56# => X"04001920",
		16#2b57# => X"15000000",
		16#2b58# => X"bc2b0000",
		16#2b59# => X"0c00015f",
		16#2b5a# => X"18800001",
		16#2b5b# => X"bc12ffff",
		16#2b5c# => X"1000023e",
		16#2b5d# => X"15000000",
		16#2b5e# => X"ae1e0047",
		16#2b5f# => X"e1608002",
		16#2b60# => X"e16b8004",
		16#2b61# => X"bd6b0000",
		16#2b62# => X"10000009",
		16#2b63# => X"bc120000",
		16#2b64# => X"ad9e0067",
		16#2b65# => X"e1606002",
		16#2b66# => X"e16b6004",
		16#2b67# => X"bd8b0000",
		16#2b68# => X"10000007",
		16#2b69# => X"84810018",
		16#2b6a# => X"bc120000",
		16#2b6b# => X"0c000004",
		16#2b6c# => X"84810018",
		16#2b6d# => X"9e400001",
		16#2b6e# => X"84810018",
		16#2b6f# => X"8441004c",
		16#2b70# => X"a8840100",
		16#2b71# => X"bd620000",
		16#2b72# => X"0c000224",
		16#2b73# => X"d4012018",
		16#2b74# => X"8701004c",
		16#2b75# => X"9f800000",
		16#2b76# => X"ac9e0046",
		16#2b77# => X"ad7e0066",
		16#2b78# => X"e0402002",
		16#2b79# => X"e0605802",
		16#2b7a# => X"e0422004",
		16#2b7b# => X"e1635804",
		16#2b7c# => X"e16b1003",
		16#2b7d# => X"ad6bffff",
		16#2b7e# => X"bb4b005f",
		16#2b7f# => X"bc3a0000",
		16#2b80# => X"100001fb",
		16#2b81# => X"a9d20000",
		16#2b82# => X"ad9e0045",
		16#2b83# => X"e1606002",
		16#2b84# => X"e16b6004",
		16#2b85# => X"bd6b0000",
		16#2b86# => X"10000009",
		16#2b87# => X"9dd20001",
		16#2b88# => X"ad9e0065",
		16#2b89# => X"e1606002",
		16#2b8a# => X"e16b6004",
		16#2b8b# => X"bd8b0000",
		16#2b8c# => X"10000211",
		16#2b8d# => X"a9d20000",
		16#2b8e# => X"9dd20001",
		16#2b8f# => X"9c400002",
		16#2b90# => X"85e10050",
		16#2b91# => X"a9980000",
		16#2b92# => X"a9af0000",
		16#2b93# => X"a8c20000",
		16#2b94# => X"9c810550",
		16#2b95# => X"84610028",
		16#2b96# => X"a8ee0000",
		16#2b97# => X"9d010554",
		16#2b98# => X"9c41054c",
		16#2b99# => X"d4012000",
		16#2b9a# => X"e08c0004",
		16#2b9b# => X"e0ad0004",
		16#2b9c# => X"0400041c",
		16#2b9d# => X"d4011004",
		16#2b9e# => X"e1a08002",
		16#2b9f# => X"e1ad8004",
		16#2ba0# => X"bd6d0000",
		16#2ba1# => X"10000008",
		16#2ba2# => X"d4015840",
		16#2ba3# => X"ad9e0067",
		16#2ba4# => X"e1a06002",
		16#2ba5# => X"e1ad6004",
		16#2ba6# => X"bd8d0000",
		16#2ba7# => X"10000007",
		16#2ba8# => X"84810040",
		16#2ba9# => X"84610018",
		16#2baa# => X"a5a30001",
		16#2bab# => X"bc2d0000",
		16#2bac# => X"0c0001f8",
		16#2bad# => X"84810040",
		16#2bae# => X"bc1a0000",
		16#2baf# => X"10000008",
		16#2bb0# => X"e0447000",
		16#2bb1# => X"91e40000",
		16#2bb2# => X"bc2f0030",
		16#2bb3# => X"0c000202",
		16#2bb4# => X"85610050",
		16#2bb5# => X"85c10554",
		16#2bb6# => X"e0427000",
		16#2bb7# => X"84810050",
		16#2bb8# => X"18600001",
		16#2bb9# => X"a9980000",
		16#2bba# => X"a8633ee4",
		16#2bbb# => X"a9a40000",
		16#2bbc# => X"84a30000",
		16#2bbd# => X"84c30004",
		16#2bbe# => X"e06c0004",
		16#2bbf# => X"e08d0004",
		16#2bc0# => X"07fff02f",
		16#2bc1# => X"15000000",
		16#2bc2# => X"bc0b0000",
		16#2bc3# => X"0c0001ba",
		16#2bc4# => X"8461054c",
		16#2bc5# => X"d401154c",
		16#2bc6# => X"a8620000",
		16#2bc7# => X"84810040",
		16#2bc8# => X"e0408002",
		16#2bc9# => X"e0632002",
		16#2bca# => X"e1028004",
		16#2bcb# => X"bd680000",
		16#2bcc# => X"10000008",
		16#2bcd# => X"d4011838",
		16#2bce# => X"ad7e0067",
		16#2bcf# => X"e1005802",
		16#2bd0# => X"e1085804",
		16#2bd1# => X"bd880000",
		16#2bd2# => X"1000019a",
		16#2bd3# => X"bc1e0066",
		16#2bd4# => X"87410554",
		16#2bd5# => X"bd9afffd",
		16#2bd6# => X"10000005",
		16#2bd7# => X"a9da0000",
		16#2bd8# => X"e572d000",
		16#2bd9# => X"1000010c",
		16#2bda# => X"84810038",
		16#2bdb# => X"9e9efffe",
		16#2bdc# => X"9dceffff",
		16#2bdd# => X"d801a544",
		16#2bde# => X"bd6e0000",
		16#2bdf# => X"0c0001cf",
		16#2be0# => X"d4017554",
		16#2be1# => X"9c60002b",
		16#2be2# => X"d8011d45",
		16#2be3# => X"bdae0009",
		16#2be4# => X"100001bb",
		16#2be5# => X"9c800030",
		16#2be6# => X"9c41046f",
		16#2be7# => X"a86e0000",
		16#2be8# => X"9c80000a",
		16#2be9# => X"04002265",
		16#2bea# => X"9c42ffff",
		16#2beb# => X"9d6b0030",
		16#2bec# => X"a86e0000",
		16#2bed# => X"9c80000a",
		16#2bee# => X"07ffe712",
		16#2bef# => X"d8025800",
		16#2bf0# => X"bd4b0009",
		16#2bf1# => X"13fffff6",
		16#2bf2# => X"a9cb0000",
		16#2bf3# => X"9d02ffff",
		16#2bf4# => X"9dcb0030",
		16#2bf5# => X"d8087000",
		16#2bf6# => X"8481000c",
		16#2bf7# => X"e4682000",
		16#2bf8# => X"10000009",
		16#2bf9# => X"9ca10546",
		16#2bfa# => X"8c480000",
		16#2bfb# => X"d8051000",
		16#2bfc# => X"9d080001",
		16#2bfd# => X"8461000c",
		16#2bfe# => X"e4881800",
		16#2bff# => X"13fffffb",
		16#2c00# => X"9ca50001",
		16#2c01# => X"84410008",
		16#2c02# => X"84610038",
		16#2c03# => X"e0a51002",
		16#2c04# => X"bd430001",
		16#2c05# => X"d4012858",
		16#2c06# => X"100000e7",
		16#2c07# => X"e3451800",
		16#2c08# => X"84810018",
		16#2c09# => X"a5040001",
		16#2c0a# => X"bc080000",
		16#2c0b# => X"0c0000e2",
		16#2c0c# => X"15000000",
		16#2c0d# => X"bc1c0000",
		16#2c0e# => X"10000144",
		16#2c0f# => X"ac5affff",
		16#2c10# => X"9c60002d",
		16#2c11# => X"b842009f",
		16#2c12# => X"9c800000",
		16#2c13# => X"d8011d5b",
		16#2c14# => X"e05a1003",
		16#2c15# => X"abd40000",
		16#2c16# => X"d4012044",
		16#2c17# => X"03fffb1a",
		16#2c18# => X"d4011024",
		16#2c19# => X"84610018",
		16#2c1a# => X"a4430040",
		16#2c1b# => X"bc020000",
		16#2c1c# => X"10000096",
		16#2c1d# => X"8481002c",
		16#2c1e# => X"84610030",
		16#2c1f# => X"84440000",
		16#2c20# => X"9c840004",
		16#2c21# => X"d401202c",
		16#2c22# => X"03fff9cb",
		16#2c23# => X"dc021800",
		16#2c24# => X"9d000001",
		16#2c25# => X"85c20000",
		16#2c26# => X"9c420004",
		16#2c27# => X"e1607002",
		16#2c28# => X"d401102c",
		16#2c29# => X"e0eb7004",
		16#2c2a# => X"03fffbbc",
		16#2c2b# => X"b967005f",
		16#2c2c# => X"a90b0000",
		16#2c2d# => X"85c30000",
		16#2c2e# => X"9c630004",
		16#2c2f# => X"e1607002",
		16#2c30# => X"d401182c",
		16#2c31# => X"e0eb7004",
		16#2c32# => X"03fffbb4",
		16#2c33# => X"b967005f",
		16#2c34# => X"a8b80000",
		16#2c35# => X"8601053c",
		16#2c36# => X"9f180008",
		16#2c37# => X"aa944050",
		16#2c38# => X"9e100001",
		16#2c39# => X"e2527000",
		16#2c3a# => X"d405a000",
		16#2c3b# => X"d4057004",
		16#2c3c# => X"d4019540",
		16#2c3d# => X"bdb00007",
		16#2c3e# => X"1000000a",
		16#2c3f# => X"d401853c",
		16#2c40# => X"84610028",
		16#2c41# => X"84810020",
		16#2c42# => X"04001934",
		16#2c43# => X"9ca10538",
		16#2c44# => X"bc2b0000",
		16#2c45# => X"13fffa5b",
		16#2c46# => X"9f0104d0",
		16#2c47# => X"86410540",
		16#2c48# => X"84410018",
		16#2c49# => X"a4a20001",
		16#2c4a# => X"bc050000",
		16#2c4b# => X"13fffc85",
		16#2c4c# => X"84810018",
		16#2c4d# => X"8601053c",
		16#2c4e# => X"84610054",
		16#2c4f# => X"9e100001",
		16#2c50# => X"e2521800",
		16#2c51# => X"84810048",
		16#2c52# => X"d4182000",
		16#2c53# => X"d4181804",
		16#2c54# => X"d4019540",
		16#2c55# => X"bd500007",
		16#2c56# => X"13fffd83",
		16#2c57# => X"d401853c",
		16#2c58# => X"03fffc77",
		16#2c59# => X"9f180008",
		16#2c5a# => X"1a800001",
		16#2c5b# => X"a8b80000",
		16#2c5c# => X"03fffc5b",
		16#2c5d# => X"aa944050",
		16#2c5e# => X"84610028",
		16#2c5f# => X"84810020",
		16#2c60# => X"04001916",
		16#2c61# => X"9ca10538",
		16#2c62# => X"bc2b0000",
		16#2c63# => X"13fffa3d",
		16#2c64# => X"9f0104d0",
		16#2c65# => X"03fffccf",
		16#2c66# => X"86410540",
		16#2c67# => X"19000001",
		16#2c68# => X"9e100001",
		16#2c69# => X"9e520001",
		16#2c6a# => X"a9083edf",
		16#2c6b# => X"9c800001",
		16#2c6c# => X"d4164000",
		16#2c6d# => X"d4162004",
		16#2c6e# => X"d4019540",
		16#2c6f# => X"bdb00007",
		16#2c70# => X"0c000060",
		16#2c71# => X"d401853c",
		16#2c72# => X"bc2e0000",
		16#2c73# => X"10000009",
		16#2c74# => X"84410038",
		16#2c75# => X"bc220000",
		16#2c76# => X"10000006",
		16#2c77# => X"84610018",
		16#2c78# => X"a5030001",
		16#2c79# => X"bc080000",
		16#2c7a# => X"13fffc56",
		16#2c7b# => X"84810018",
		16#2c7c# => X"8601053c",
		16#2c7d# => X"84810054",
		16#2c7e# => X"9e100001",
		16#2c7f# => X"e2522000",
		16#2c80# => X"84410048",
		16#2c81# => X"d4182004",
		16#2c82# => X"d4181000",
		16#2c83# => X"d4019540",
		16#2c84# => X"bd500007",
		16#2c85# => X"10000055",
		16#2c86# => X"d401853c",
		16#2c87# => X"9f180008",
		16#2c88# => X"e1c07002",
		16#2c89# => X"bdae0000",
		16#2c8a# => X"1000007c",
		16#2c8b# => X"bdae0010",
		16#2c8c# => X"10000094",
		16#2c8d# => X"1a800001",
		16#2c8e# => X"9c400010",
		16#2c8f# => X"aa944050",
		16#2c90# => X"86c10028",
		16#2c91# => X"00000007",
		16#2c92# => X"87410020",
		16#2c93# => X"9f180008",
		16#2c94# => X"9dcefff0",
		16#2c95# => X"bd4e0010",
		16#2c96# => X"0c00008b",
		16#2c97# => X"15000000",
		16#2c98# => X"9e100001",
		16#2c99# => X"9e520010",
		16#2c9a# => X"d418a000",
		16#2c9b# => X"d4181004",
		16#2c9c# => X"d4019540",
		16#2c9d# => X"bd500007",
		16#2c9e# => X"0ffffff5",
		16#2c9f# => X"d401853c",
		16#2ca0# => X"a8760000",
		16#2ca1# => X"a89a0000",
		16#2ca2# => X"040018d4",
		16#2ca3# => X"9ca10538",
		16#2ca4# => X"bc2b0000",
		16#2ca5# => X"13fff9fb",
		16#2ca6# => X"9f0104d0",
		16#2ca7# => X"86410540",
		16#2ca8# => X"03ffffec",
		16#2ca9# => X"8601053c",
		16#2caa# => X"9c800000",
		16#2cab# => X"b842009f",
		16#2cac# => X"9101055b",
		16#2cad# => X"e05a1003",
		16#2cae# => X"d401702c",
		16#2caf# => X"d4012044",
		16#2cb0# => X"03fffa7e",
		16#2cb1# => X"d4011024",
		16#2cb2# => X"84610030",
		16#2cb3# => X"84440000",
		16#2cb4# => X"9c840004",
		16#2cb5# => X"d401202c",
		16#2cb6# => X"03fff937",
		16#2cb7# => X"d4021800",
		16#2cb8# => X"bd5e0047",
		16#2cb9# => X"a8843eb2",
		16#2cba# => X"10000005",
		16#2cbb# => X"d4012040",
		16#2cbc# => X"18400001",
		16#2cbd# => X"a8423eae",
		16#2cbe# => X"d4011040",
		16#2cbf# => X"9c600003",
		16#2cc0# => X"84810018",
		16#2cc1# => X"9c40ff7f",
		16#2cc2# => X"d4011824",
		16#2cc3# => X"e0841003",
		16#2cc4# => X"ab430000",
		16#2cc5# => X"9c600000",
		16#2cc6# => X"d4012018",
		16#2cc7# => X"9101055b",
		16#2cc8# => X"03fffa66",
		16#2cc9# => X"d4011844",
		16#2cca# => X"9d00002d",
		16#2ccb# => X"03fffa90",
		16#2ccc# => X"d8011d5b",
		16#2ccd# => X"ab580000",
		16#2cce# => X"03fffd49",
		16#2ccf# => X"9f180008",
		16#2cd0# => X"84610028",
		16#2cd1# => X"84810020",
		16#2cd2# => X"040018a4",
		16#2cd3# => X"9ca10538",
		16#2cd4# => X"bc2b0000",
		16#2cd5# => X"13fff9cb",
		16#2cd6# => X"85c10554",
		16#2cd7# => X"9f0104d0",
		16#2cd8# => X"03ffff9a",
		16#2cd9# => X"86410540",
		16#2cda# => X"84610028",
		16#2cdb# => X"84810020",
		16#2cdc# => X"0400189a",
		16#2cdd# => X"9ca10538",
		16#2cde# => X"bc2b0000",
		16#2cdf# => X"13fff9c1",
		16#2ce0# => X"85c10554",
		16#2ce1# => X"9f0104d0",
		16#2ce2# => X"86410540",
		16#2ce3# => X"03ffffa5",
		16#2ce4# => X"8601053c",
		16#2ce5# => X"e59a2000",
		16#2ce6# => X"100000c0",
		16#2ce7# => X"bd4e0000",
		16#2ce8# => X"84610018",
		16#2ce9# => X"a4430001",
		16#2cea# => X"bc020000",
		16#2ceb# => X"13ffff22",
		16#2cec# => X"9e800067",
		16#2ced# => X"03ffff20",
		16#2cee# => X"9f5a0001",
		16#2cef# => X"9f0e0008",
		16#2cf0# => X"03fffd27",
		16#2cf1# => X"ab4e0000",
		16#2cf2# => X"84610028",
		16#2cf3# => X"84810020",
		16#2cf4# => X"04001882",
		16#2cf5# => X"9ca10538",
		16#2cf6# => X"bc2b0000",
		16#2cf7# => X"13fff9a9",
		16#2cf8# => X"86410540",
		16#2cf9# => X"03fffc50",
		16#2cfa# => X"9ca104d0",
		16#2cfb# => X"03fffbd4",
		16#2cfc# => X"ab050000",
		16#2cfd# => X"84610028",
		16#2cfe# => X"84810020",
		16#2cff# => X"04001877",
		16#2d00# => X"9ca10538",
		16#2d01# => X"bc2b0000",
		16#2d02# => X"13fff99e",
		16#2d03# => X"9f0104d0",
		16#2d04# => X"86410540",
		16#2d05# => X"8601053c",
		16#2d06# => X"84610038",
		16#2d07# => X"9e100001",
		16#2d08# => X"e2521800",
		16#2d09# => X"03ffff49",
		16#2d0a# => X"84810040",
		16#2d0b# => X"07fff852",
		16#2d0c# => X"d401702c",
		16#2d0d# => X"adabffff",
		16#2d0e# => X"9c400000",
		16#2d0f# => X"b9ad009f",
		16#2d10# => X"ab4b0000",
		16#2d11# => X"9101055b",
		16#2d12# => X"e1ab6803",
		16#2d13# => X"d4011044",
		16#2d14# => X"03fffa1a",
		16#2d15# => X"d4016824",
		16#2d16# => X"1a800001",
		16#2d17# => X"9cf60008",
		16#2d18# => X"86410540",
		16#2d19# => X"8601053c",
		16#2d1a# => X"03fff956",
		16#2d1b# => X"aa944060",
		16#2d1c# => X"84610014",
		16#2d1d# => X"84810040",
		16#2d1e# => X"03fffa0a",
		16#2d1f# => X"e3432002",
		16#2d20# => X"aa944050",
		16#2d21# => X"9e100001",
		16#2d22# => X"e2527000",
		16#2d23# => X"d418a000",
		16#2d24# => X"d4187004",
		16#2d25# => X"d4019540",
		16#2d26# => X"bd500007",
		16#2d27# => X"13ffffd6",
		16#2d28# => X"d401853c",
		16#2d29# => X"03ffffdd",
		16#2d2a# => X"9f180008",
		16#2d2b# => X"bcb20006",
		16#2d2c# => X"10000003",
		16#2d2d# => X"ab520000",
		16#2d2e# => X"9f400006",
		16#2d2f# => X"ac5affff",
		16#2d30# => X"18800001",
		16#2d31# => X"b842009f",
		16#2d32# => X"a8843ed8",
		16#2d33# => X"d401702c",
		16#2d34# => X"e05a1003",
		16#2d35# => X"d4012040",
		16#2d36# => X"03fff8fd",
		16#2d37# => X"d4011024",
		16#2d38# => X"84610028",
		16#2d39# => X"9c40ffff",
		16#2d3a# => X"040000ac",
		16#2d3b# => X"d4011030",
		16#2d3c# => X"bc2b0000",
		16#2d3d# => X"13fff96b",
		16#2d3e# => X"84610020",
		16#2d3f# => X"9843000c",
		16#2d40# => X"03fff88f",
		16#2d41# => X"a4e2ffff",
		16#2d42# => X"1a800001",
		16#2d43# => X"8601053c",
		16#2d44# => X"03fffbb7",
		16#2d45# => X"aa944060",
		16#2d46# => X"84610028",
		16#2d47# => X"84810020",
		16#2d48# => X"0400182e",
		16#2d49# => X"9ca10538",
		16#2d4a# => X"bc2b0000",
		16#2d4b# => X"13fff955",
		16#2d4c# => X"85c10554",
		16#2d4d# => X"85610540",
		16#2d4e# => X"a84e0000",
		16#2d4f# => X"8601053c",
		16#2d50# => X"03fffc70",
		16#2d51# => X"9f0104d0",
		16#2d52# => X"9101055b",
		16#2d53# => X"b842009f",
		16#2d54# => X"abd40000",
		16#2d55# => X"d401e044",
		16#2d56# => X"e05a1003",
		16#2d57# => X"03fff9d7",
		16#2d58# => X"d4011024",
		16#2d59# => X"84610028",
		16#2d5a# => X"84810020",
		16#2d5b# => X"0400181b",
		16#2d5c# => X"9ca10538",
		16#2d5d# => X"bc2b0000",
		16#2d5e# => X"13fff942",
		16#2d5f# => X"85c10554",
		16#2d60# => X"03fffc6b",
		16#2d61# => X"9f0104d0",
		16#2d62# => X"84610028",
		16#2d63# => X"84810020",
		16#2d64# => X"04001812",
		16#2d65# => X"9ca10538",
		16#2d66# => X"bc2b0000",
		16#2d67# => X"13fff939",
		16#2d68# => X"85c10554",
		16#2d69# => X"9f0104d0",
		16#2d6a# => X"03fffd04",
		16#2d6b# => X"86410540",
		16#2d6c# => X"0c000046",
		16#2d6d# => X"15000000",
		16#2d6e# => X"87410554",
		16#2d6f# => X"bdba0000",
		16#2d70# => X"1000005c",
		16#2d71# => X"bc320000",
		16#2d72# => X"10000006",
		16#2d73# => X"84410018",
		16#2d74# => X"a5020001",
		16#2d75# => X"bc080000",
		16#2d76# => X"13fffe98",
		16#2d77# => X"bc1c0000",
		16#2d78# => X"9f5a0001",
		16#2d79# => X"03fffe94",
		16#2d7a# => X"e35a9000",
		16#2d7b# => X"03fffe15",
		16#2d7c# => X"9c400003",
		16#2d7d# => X"e4a21800",
		16#2d7e# => X"13fffe49",
		16#2d7f# => X"a8e30000",
		16#2d80# => X"9c800030",
		16#2d81# => X"d8072000",
		16#2d82# => X"9ce70001",
		16#2d83# => X"e4423800",
		16#2d84# => X"13fffffd",
		16#2d85# => X"d4013d4c",
		16#2d86# => X"9da30001",
		16#2d87# => X"9c800001",
		16#2d88# => X"e1a46802",
		16#2d89# => X"e1a26800",
		16#2d8a# => X"03fffe3d",
		16#2d8b# => X"e0636800",
		16#2d8c# => X"1a800001",
		16#2d8d# => X"a9180000",
		16#2d8e# => X"03fffc15",
		16#2d8f# => X"aa944050",
		16#2d90# => X"d4019024",
		16#2d91# => X"9101055b",
		16#2d92# => X"ab520000",
		16#2d93# => X"d401702c",
		16#2d94# => X"03fff99a",
		16#2d95# => X"d4015844",
		16#2d96# => X"18608000",
		16#2d97# => X"9f80002d",
		16#2d98# => X"03fffdde",
		16#2d99# => X"e3021800",
		16#2d9a# => X"9e400006",
		16#2d9b# => X"03fffdd3",
		16#2d9c# => X"ae1e0047",
		16#2d9d# => X"03fffdf3",
		16#2d9e# => X"9c400002",
		16#2d9f# => X"9dce0030",
		16#2da0# => X"d8017547",
		16#2da1# => X"d8012546",
		16#2da2# => X"03fffe5f",
		16#2da3# => X"9ca10548",
		16#2da4# => X"03fffe23",
		16#2da5# => X"8461054c",
		16#2da6# => X"10000004",
		16#2da7# => X"9f400001",
		16#2da8# => X"9c800002",
		16#2da9# => X"e3447002",
		16#2daa# => X"84410038",
		16#2dab# => X"9e800067",
		16#2dac# => X"03fffe61",
		16#2dad# => X"e35a1000",
		16#2dae# => X"9c40002d",
		16#2daf# => X"e1c07002",
		16#2db0# => X"03fffe33",
		16#2db1# => X"d8011545",
		16#2db2# => X"aa9e0000",
		16#2db3# => X"03fffe29",
		16#2db4# => X"85c10554",
		16#2db5# => X"18600001",
		16#2db6# => X"a9980000",
		16#2db7# => X"a8633ee4",
		16#2db8# => X"a9ab0000",
		16#2db9# => X"84a30000",
		16#2dba# => X"84c30004",
		16#2dbb# => X"e06c0004",
		16#2dbc# => X"e08d0004",
		16#2dbd# => X"07ffee50",
		16#2dbe# => X"15000000",
		16#2dbf# => X"bc2b0000",
		16#2dc0# => X"0ffffdf5",
		16#2dc1# => X"9c800001",
		16#2dc2# => X"e1c47002",
		16#2dc3# => X"03fffdf2",
		16#2dc4# => X"d4017554",
		16#2dc5# => X"8441002c",
		16#2dc6# => X"86420000",
		16#2dc7# => X"bd920000",
		16#2dc8# => X"1000000f",
		16#2dc9# => X"9c420004",
		16#2dca# => X"03fff857",
		16#2dcb# => X"d401102c",
		16#2dcc# => X"13fffe41",
		16#2dcd# => X"9f520002",
		16#2dce# => X"84610018",
		16#2dcf# => X"a4430001",
		16#2dd0# => X"bc020000",
		16#2dd1# => X"13fffe3c",
		16#2dd2# => X"9f400001",
		16#2dd3# => X"03fffe3a",
		16#2dd4# => X"9f520002",
		16#2dd5# => X"03fff905",
		16#2dd6# => X"d4011830",
		16#2dd7# => X"d401102c",
		16#2dd8# => X"03fff849",
		16#2dd9# => X"9e40ffff",
		16#2dda# => X"a8e40000",
		16#2ddb# => X"a8830000",
		16#2ddc# => X"18600001",
		16#2ddd# => X"d7e14ffc",
		16#2dde# => X"a86363e0",
		16#2ddf# => X"9c21fffc",
		16#2de0# => X"84630000",
		16#2de1# => X"9c210004",
		16#2de2# => X"a8c50000",
		16#2de3# => X"8521fffc",
		16#2de4# => X"03fff7b7",
		16#2de5# => X"a8a70000",
		16#2de6# => X"d7e117f4",
		16#2de7# => X"18400001",
		16#2de8# => X"d7e177f8",
		16#2de9# => X"a84263e0",
		16#2dea# => X"d7e14ffc",
		16#2deb# => X"84a20000",
		16#2dec# => X"9c21fff4",
		16#2ded# => X"a9c30000",
		16#2dee# => X"bc050000",
		16#2def# => X"10000006",
		16#2df0# => X"a8440000",
		16#2df1# => X"84650038",
		16#2df2# => X"bc230000",
		16#2df3# => X"0c00002b",
		16#2df4# => X"15000000",
		16#2df5# => X"98c2000c",
		16#2df6# => X"a486ffff",
		16#2df7# => X"a4640008",
		16#2df8# => X"bc030000",
		16#2df9# => X"10000032",
		16#2dfa# => X"a8e60000",
		16#2dfb# => X"84a20010",
		16#2dfc# => X"bc250000",
		16#2dfd# => X"0c000025",
		16#2dfe# => X"a4640280",
		16#2dff# => X"a4640001",
		16#2e00# => X"bc030000",
		16#2e01# => X"1000000f",
		16#2e02# => X"a4840002",
		16#2e03# => X"84620014",
		16#2e04# => X"9c800000",
		16#2e05# => X"e0601802",
		16#2e06# => X"9d600000",
		16#2e07# => X"d4022008",
		16#2e08# => X"e4255800",
		16#2e09# => X"0c00000e",
		16#2e0a# => X"d4021818",
		16#2e0b# => X"9c21000c",
		16#2e0c# => X"8521fffc",
		16#2e0d# => X"8441fff4",
		16#2e0e# => X"44004800",
		16#2e0f# => X"85c1fff8",
		16#2e10# => X"bc240000",
		16#2e11# => X"10000003",
		16#2e12# => X"9d600000",
		16#2e13# => X"84620014",
		16#2e14# => X"e4255800",
		16#2e15# => X"13fffff6",
		16#2e16# => X"d4021808",
		16#2e17# => X"9442000c",
		16#2e18# => X"a4420080",
		16#2e19# => X"bc220000",
		16#2e1a# => X"13fffff1",
		16#2e1b# => X"9d60ffff",
		16#2e1c# => X"03ffffef",
		16#2e1d# => X"a9650000",
		16#2e1e# => X"040009d0",
		16#2e1f# => X"a8650000",
		16#2e20# => X"03ffffd6",
		16#2e21# => X"98c2000c",
		16#2e22# => X"bc030200",
		16#2e23# => X"13ffffdd",
		16#2e24# => X"a4640001",
		16#2e25# => X"a8820000",
		16#2e26# => X"04000dcb",
		16#2e27# => X"a86e0000",
		16#2e28# => X"9482000c",
		16#2e29# => X"03ffffd6",
		16#2e2a# => X"84a20010",
		16#2e2b# => X"a4640010",
		16#2e2c# => X"bc030000",
		16#2e2d# => X"13ffffde",
		16#2e2e# => X"9d60ffff",
		16#2e2f# => X"a4840004",
		16#2e30# => X"bc240000",
		16#2e31# => X"10000007",
		16#2e32# => X"15000000",
		16#2e33# => X"84a20010",
		16#2e34# => X"a8860008",
		16#2e35# => X"dc02200c",
		16#2e36# => X"03ffffc6",
		16#2e37# => X"a484ffff",
		16#2e38# => X"84820030",
		16#2e39# => X"bc040000",
		16#2e3a# => X"1000000a",
		16#2e3b# => X"9c620040",
		16#2e3c# => X"e4041800",
		16#2e3d# => X"10000006",
		16#2e3e# => X"9c600000",
		16#2e3f# => X"04000ad0",
		16#2e40# => X"a86e0000",
		16#2e41# => X"98e2000c",
		16#2e42# => X"9c600000",
		16#2e43# => X"d4021830",
		16#2e44# => X"84a20010",
		16#2e45# => X"9c80ffdb",
		16#2e46# => X"9c600000",
		16#2e47# => X"e0c72003",
		16#2e48# => X"d4021804",
		16#2e49# => X"03ffffeb",
		16#2e4a# => X"d4022800",
		16#2e4b# => X"d7e117e4",
		16#2e4c# => X"a8430000",
		16#2e4d# => X"18600001",
		16#2e4e# => X"d7e1b7f8",
		16#2e4f# => X"a8633ea0",
		16#2e50# => X"d7e187ec",
		16#2e51# => X"86c30000",
		16#2e52# => X"d7e197f0",
		16#2e53# => X"d7e1a7f4",
		16#2e54# => X"d7e14ffc",
		16#2e55# => X"d7e177e8",
		16#2e56# => X"84f60148",
		16#2e57# => X"9c21ffe4",
		16#2e58# => X"aa040000",
		16#2e59# => X"aa850000",
		16#2e5a# => X"bc270000",
		16#2e5b# => X"0c00002c",
		16#2e5c# => X"aa460000",
		16#2e5d# => X"85070004",
		16#2e5e# => X"bda8001f",
		16#2e5f# => X"0c00002b",
		16#2e60# => X"18600000",
		16#2e61# => X"bc020000",
		16#2e62# => X"0c000013",
		16#2e63# => X"9c880042",
		16#2e64# => X"9c480002",
		16#2e65# => X"9d080001",
		16#2e66# => X"b8420002",
		16#2e67# => X"d4074004",
		16#2e68# => X"9dc00000",
		16#2e69# => X"e0e71000",
		16#2e6a# => X"d4078000",
		16#2e6b# => X"9c21001c",
		16#2e6c# => X"a96e0000",
		16#2e6d# => X"8521fffc",
		16#2e6e# => X"8441ffe4",
		16#2e6f# => X"85c1ffe8",
		16#2e70# => X"8601ffec",
		16#2e71# => X"8641fff0",
		16#2e72# => X"8681fff4",
		16#2e73# => X"44004800",
		16#2e74# => X"86c1fff8",
		16#2e75# => X"9cc80022",
		16#2e76# => X"9c600001",
		16#2e77# => X"b8c60002",
		16#2e78# => X"e0634008",
		16#2e79# => X"b8840002",
		16#2e7a# => X"84a70188",
		16#2e7b# => X"e0c73000",
		16#2e7c# => X"e0a51804",
		16#2e7d# => X"e0872000",
		16#2e7e# => X"d406a000",
		16#2e7f# => X"d4072988",
		16#2e80# => X"bc220002",
		16#2e81# => X"13ffffe3",
		16#2e82# => X"d4049000",
		16#2e83# => X"8447018c",
		16#2e84# => X"e0621804",
		16#2e85# => X"03ffffdf",
		16#2e86# => X"d407198c",
		16#2e87# => X"9cf6014c",
		16#2e88# => X"03ffffd5",
		16#2e89# => X"d4163948",
		16#2e8a# => X"a8637918",
		16#2e8b# => X"bc030000",
		16#2e8c# => X"13ffffdf",
		16#2e8d# => X"9dc0ffff",
		16#2e8e# => X"07ffefb8",
		16#2e8f# => X"9c600190",
		16#2e90# => X"bc0b0000",
		16#2e91# => X"13ffffda",
		16#2e92# => X"a8eb0000",
		16#2e93# => X"84760148",
		16#2e94# => X"9c800000",
		16#2e95# => X"d40b1800",
		16#2e96# => X"d40b2004",
		16#2e97# => X"d4165948",
		16#2e98# => X"d40b2188",
		16#2e99# => X"d40b218c",
		16#2e9a# => X"03ffffc7",
		16#2e9b# => X"a9040000",
		16#2e9c# => X"d7e117d4",
		16#2e9d# => X"18400001",
		16#2e9e# => X"d7e1f7f8",
		16#2e9f# => X"a8423ea0",
		16#2ea0# => X"d7e1a7e4",
		16#2ea1# => X"87c20000",
		16#2ea2# => X"d7e1d7f0",
		16#2ea3# => X"d7e1e7f4",
		16#2ea4# => X"d7e14ffc",
		16#2ea5# => X"d7e177d8",
		16#2ea6# => X"d7e187dc",
		16#2ea7# => X"d7e197e0",
		16#2ea8# => X"d7e1b7e8",
		16#2ea9# => X"d7e1c7ec",
		16#2eaa# => X"9c5e0148",
		16#2eab# => X"9c21ffd0",
		16#2eac# => X"ab830000",
		16#2ead# => X"aa840000",
		16#2eae# => X"d4011000",
		16#2eaf# => X"9f400001",
		16#2eb0# => X"85de0148",
		16#2eb1# => X"bc0e0000",
		16#2eb2# => X"10000041",
		16#2eb3# => X"86c10000",
		16#2eb4# => X"848e0004",
		16#2eb5# => X"9c44ffff",
		16#2eb6# => X"bd820000",
		16#2eb7# => X"10000037",
		16#2eb8# => X"15000000",
		16#2eb9# => X"9e040021",
		16#2eba# => X"9e440001",
		16#2ebb# => X"ba100002",
		16#2ebc# => X"ba520002",
		16#2ebd# => X"e20e8000",
		16#2ebe# => X"0000000b",
		16#2ebf# => X"e24e9000",
		16#2ec0# => X"84900080",
		16#2ec1# => X"e424a000",
		16#2ec2# => X"0c00000a",
		16#2ec3# => X"15000000",
		16#2ec4# => X"9c42ffff",
		16#2ec5# => X"9e10fffc",
		16#2ec6# => X"bd620000",
		16#2ec7# => X"0c000027",
		16#2ec8# => X"9e52fffc",
		16#2ec9# => X"bc140000",
		16#2eca# => X"0ffffff6",
		16#2ecb# => X"15000000",
		16#2ecc# => X"848e0004",
		16#2ecd# => X"9c84ffff",
		16#2ece# => X"e4241000",
		16#2ecf# => X"0c000035",
		16#2ed0# => X"84b20000",
		16#2ed1# => X"9c600000",
		16#2ed2# => X"d4121800",
		16#2ed3# => X"bc050000",
		16#2ed4# => X"13fffff0",
		16#2ed5# => X"e09a1008",
		16#2ed6# => X"84ce0188",
		16#2ed7# => X"e0c43003",
		16#2ed8# => X"bc260000",
		16#2ed9# => X"0c000027",
		16#2eda# => X"870e0004",
		16#2edb# => X"84ce018c",
		16#2edc# => X"e0843003",
		16#2edd# => X"bc240000",
		16#2ede# => X"10000028",
		16#2edf# => X"a87c0000",
		16#2ee0# => X"48002800",
		16#2ee1# => X"84900000",
		16#2ee2# => X"848e0004",
		16#2ee3# => X"e424c000",
		16#2ee4# => X"13ffffcc",
		16#2ee5# => X"15000000",
		16#2ee6# => X"84960000",
		16#2ee7# => X"e4247000",
		16#2ee8# => X"13ffffc8",
		16#2ee9# => X"9c42ffff",
		16#2eea# => X"9e10fffc",
		16#2eeb# => X"bd620000",
		16#2eec# => X"13ffffdd",
		16#2eed# => X"9e52fffc",
		16#2eee# => X"18400000",
		16#2eef# => X"a8427940",
		16#2ef0# => X"bc020000",
		16#2ef1# => X"0c000019",
		16#2ef2# => X"15000000",
		16#2ef3# => X"9c210030",
		16#2ef4# => X"8521fffc",
		16#2ef5# => X"8441ffd4",
		16#2ef6# => X"85c1ffd8",
		16#2ef7# => X"8601ffdc",
		16#2ef8# => X"8641ffe0",
		16#2ef9# => X"8681ffe4",
		16#2efa# => X"86c1ffe8",
		16#2efb# => X"8701ffec",
		16#2efc# => X"8741fff0",
		16#2efd# => X"8781fff4",
		16#2efe# => X"44004800",
		16#2eff# => X"87c1fff8",
		16#2f00# => X"48002800",
		16#2f01# => X"15000000",
		16#2f02# => X"03ffffe1",
		16#2f03# => X"848e0004",
		16#2f04# => X"03ffffcf",
		16#2f05# => X"d40e1004",
		16#2f06# => X"48002800",
		16#2f07# => X"84700000",
		16#2f08# => X"03ffffdb",
		16#2f09# => X"848e0004",
		16#2f0a# => X"844e0004",
		16#2f0b# => X"bc220000",
		16#2f0c# => X"0c00000a",
		16#2f0d# => X"15000000",
		16#2f0e# => X"844e0000",
		16#2f0f# => X"aace0000",
		16#2f10# => X"a9c20000",
		16#2f11# => X"bc2e0000",
		16#2f12# => X"13ffffa2",
		16#2f13# => X"15000000",
		16#2f14# => X"03ffffe0",
		16#2f15# => X"9c210030",
		16#2f16# => X"844e0000",
		16#2f17# => X"bc020000",
		16#2f18# => X"13fffff7",
		16#2f19# => X"a86e0000",
		16#2f1a# => X"07ffef36",
		16#2f1b# => X"d4161000",
		16#2f1c# => X"03fffff5",
		16#2f1d# => X"85d60000",
		16#2f1e# => X"d7e117dc",
		16#2f1f# => X"d7e177e0",
		16#2f20# => X"d7e187e4",
		16#2f21# => X"d7e1b7f0",
		16#2f22# => X"d7e1d7f8",
		16#2f23# => X"d7e14ffc",
		16#2f24# => X"d7e197e8",
		16#2f25# => X"d7e1a7ec",
		16#2f26# => X"d7e1c7f4",
		16#2f27# => X"84430010",
		16#2f28# => X"85c40010",
		16#2f29# => X"9c21ffdc",
		16#2f2a# => X"aa030000",
		16#2f2b# => X"aac40000",
		16#2f2c# => X"e54e1000",
		16#2f2d# => X"1000007f",
		16#2f2e# => X"9f400000",
		16#2f2f# => X"9c6e0004",
		16#2f30# => X"9c440014",
		16#2f31# => X"b8630002",
		16#2f32# => X"9dceffff",
		16#2f33# => X"9f100014",
		16#2f34# => X"e2441800",
		16#2f35# => X"e0701800",
		16#2f36# => X"84920000",
		16#2f37# => X"84630000",
		16#2f38# => X"07ffe389",
		16#2f39# => X"9c840001",
		16#2f3a# => X"e40bd000",
		16#2f3b# => X"1000003b",
		16#2f3c# => X"aa8b0000",
		16#2f3d# => X"a97a0000",
		16#2f3e# => X"a8c20000",
		16#2f3f# => X"a8b80000",
		16#2f40# => X"a87a0000",
		16#2f41# => X"85860000",
		16#2f42# => X"85050000",
		16#2f43# => X"a4ecffff",
		16#2f44# => X"b98c0050",
		16#2f45# => X"e0f43b06",
		16#2f46# => X"e1946306",
		16#2f47# => X"e0eb3800",
		16#2f48# => X"a488ffff",
		16#2f49# => X"b9670050",
		16#2f4a# => X"e0632000",
		16#2f4b# => X"a4e7ffff",
		16#2f4c# => X"e16b6000",
		16#2f4d# => X"e0833802",
		16#2f4e# => X"b8680050",
		16#2f4f# => X"a50bffff",
		16#2f50# => X"b8e40090",
		16#2f51# => X"e0634002",
		16#2f52# => X"a484ffff",
		16#2f53# => X"e0633800",
		16#2f54# => X"9cc60004",
		16#2f55# => X"b8e30010",
		16#2f56# => X"b96b0050",
		16#2f57# => X"b8630090",
		16#2f58# => X"e0872004",
		16#2f59# => X"e4723000",
		16#2f5a# => X"d4052000",
		16#2f5b# => X"13ffffe6",
		16#2f5c# => X"9ca50004",
		16#2f5d# => X"9cae0005",
		16#2f5e# => X"b8a50002",
		16#2f5f# => X"e0b02800",
		16#2f60# => X"84650000",
		16#2f61# => X"bc230000",
		16#2f62# => X"10000015",
		16#2f63# => X"a8700000",
		16#2f64# => X"9ca5fffc",
		16#2f65# => X"e4782800",
		16#2f66# => X"1000000f",
		16#2f67# => X"15000000",
		16#2f68# => X"84650000",
		16#2f69# => X"bc230000",
		16#2f6a# => X"0c000008",
		16#2f6b# => X"9ca5fffc",
		16#2f6c# => X"0000000a",
		16#2f6d# => X"d4107010",
		16#2f6e# => X"84650000",
		16#2f6f# => X"bc030000",
		16#2f70# => X"0c000005",
		16#2f71# => X"9ca5fffc",
		16#2f72# => X"e4782800",
		16#2f73# => X"0ffffffb",
		16#2f74# => X"9dceffff",
		16#2f75# => X"d4107010",
		16#2f76# => X"a8700000",
		16#2f77# => X"040010b4",
		16#2f78# => X"a8960000",
		16#2f79# => X"bd8b0000",
		16#2f7a# => X"10000031",
		16#2f7b# => X"a8980000",
		16#2f7c# => X"9e940001",
		16#2f7d# => X"9c600000",
		16#2f7e# => X"84e20000",
		16#2f7f# => X"85040000",
		16#2f80# => X"a4a7ffff",
		16#2f81# => X"a4c8ffff",
		16#2f82# => X"b8e70050",
		16#2f83# => X"e0a62802",
		16#2f84# => X"b9080050",
		16#2f85# => X"e0a51800",
		16#2f86# => X"9c420004",
		16#2f87# => X"b8c50090",
		16#2f88# => X"e0683802",
		16#2f89# => X"a4a5ffff",
		16#2f8a# => X"e0633000",
		16#2f8b# => X"e4721000",
		16#2f8c# => X"b8c30010",
		16#2f8d# => X"b8630090",
		16#2f8e# => X"e0a62804",
		16#2f8f# => X"d4042800",
		16#2f90# => X"13ffffee",
		16#2f91# => X"9c840004",
		16#2f92# => X"9c4e0005",
		16#2f93# => X"b8420002",
		16#2f94# => X"e0501000",
		16#2f95# => X"84620000",
		16#2f96# => X"bc230000",
		16#2f97# => X"10000015",
		16#2f98# => X"ab540000",
		16#2f99# => X"9c42fffc",
		16#2f9a# => X"e4781000",
		16#2f9b# => X"1000000f",
		16#2f9c# => X"15000000",
		16#2f9d# => X"84620000",
		16#2f9e# => X"bc230000",
		16#2f9f# => X"0c000008",
		16#2fa0# => X"9c42fffc",
		16#2fa1# => X"0000000b",
		16#2fa2# => X"d4107010",
		16#2fa3# => X"84620000",
		16#2fa4# => X"bc030000",
		16#2fa5# => X"0c000005",
		16#2fa6# => X"9c42fffc",
		16#2fa7# => X"e4781000",
		16#2fa8# => X"0ffffffb",
		16#2fa9# => X"9dceffff",
		16#2faa# => X"d4107010",
		16#2fab# => X"ab540000",
		16#2fac# => X"9c210024",
		16#2fad# => X"a97a0000",
		16#2fae# => X"8521fffc",
		16#2faf# => X"8441ffdc",
		16#2fb0# => X"85c1ffe0",
		16#2fb1# => X"8601ffe4",
		16#2fb2# => X"8641ffe8",
		16#2fb3# => X"8681ffec",
		16#2fb4# => X"86c1fff0",
		16#2fb5# => X"8701fff4",
		16#2fb6# => X"44004800",
		16#2fb7# => X"8741fff8",
		16#2fb8# => X"d7e117d4",
		16#2fb9# => X"d7e177d8",
		16#2fba# => X"d7e1e7f4",
		16#2fbb# => X"d7e1f7f8",
		16#2fbc# => X"d7e14ffc",
		16#2fbd# => X"d7e187dc",
		16#2fbe# => X"d7e197e0",
		16#2fbf# => X"d7e1a7e4",
		16#2fc0# => X"d7e1b7e8",
		16#2fc1# => X"d7e1c7ec",
		16#2fc2# => X"d7e1d7f0",
		16#2fc3# => X"9c21ff64",
		16#2fc4# => X"84430040",
		16#2fc5# => X"d4013000",
		16#2fc6# => X"d4013818",
		16#2fc7# => X"d4014014",
		16#2fc8# => X"d4012810",
		16#2fc9# => X"abc30000",
		16#2fca# => X"85c1009c",
		16#2fcb# => X"bc020000",
		16#2fcc# => X"1000000b",
		16#2fcd# => X"ab840000",
		16#2fce# => X"85630044",
		16#2fcf# => X"9d800001",
		16#2fd0# => X"d4025804",
		16#2fd1# => X"e16c5808",
		16#2fd2# => X"a8820000",
		16#2fd3# => X"d4025808",
		16#2fd4# => X"04000e02",
		16#2fd5# => X"9c400000",
		16#2fd6# => X"d41e1040",
		16#2fd7# => X"bd7c0000",
		16#2fd8# => X"0c000204",
		16#2fd9# => X"9c800000",
		16#2fda# => X"d40e2000",
		16#2fdb# => X"18c07ff0",
		16#2fdc# => X"e05c3003",
		16#2fdd# => X"e4223000",
		16#2fde# => X"0c0001e2",
		16#2fdf# => X"85810010",
		16#2fe0# => X"18e00001",
		16#2fe1# => X"a85c0000",
		16#2fe2# => X"a86c0000",
		16#2fe3# => X"a8e74080",
		16#2fe4# => X"e0830004",
		16#2fe5# => X"e0620004",
		16#2fe6# => X"a9cc0000",
		16#2fe7# => X"84a70000",
		16#2fe8# => X"84c70004",
		16#2fe9# => X"07ffec24",
		16#2fea# => X"aa1c0000",
		16#2feb# => X"bc2b0000",
		16#2fec# => X"0c00001d",
		16#2fed# => X"9c400001",
		16#2fee# => X"a44200ff",
		16#2fef# => X"bc220000",
		16#2ff0# => X"1000001f",
		16#2ff1# => X"ba5c0054",
		16#2ff2# => X"9c400001",
		16#2ff3# => X"84610014",
		16#2ff4# => X"19600001",
		16#2ff5# => X"848100a0",
		16#2ff6# => X"d4031000",
		16#2ff7# => X"bc040000",
		16#2ff8# => X"10000004",
		16#2ff9# => X"a96b3edf",
		16#2ffa# => X"e04b1000",
		16#2ffb# => X"d4041000",
		16#2ffc# => X"9c21009c",
		16#2ffd# => X"8521fffc",
		16#2ffe# => X"8441ffd4",
		16#2fff# => X"85c1ffd8",
		16#3000# => X"8601ffdc",
		16#3001# => X"8641ffe0",
		16#3002# => X"8681ffe4",
		16#3003# => X"86c1ffe8",
		16#3004# => X"8701ffec",
		16#3005# => X"8741fff0",
		16#3006# => X"8781fff4",
		16#3007# => X"44004800",
		16#3008# => X"87c1fff8",
		16#3009# => X"9c400000",
		16#300a# => X"a44200ff",
		16#300b# => X"bc220000",
		16#300c# => X"0fffffe7",
		16#300d# => X"9c400001",
		16#300e# => X"ba5c0054",
		16#300f# => X"a9700000",
		16#3010# => X"a98e0000",
		16#3011# => X"a87e0000",
		16#3012# => X"9cc10068",
		16#3013# => X"9ce1006c",
		16#3014# => X"e08b0004",
		16#3015# => X"e0ac0004",
		16#3016# => X"04001113",
		16#3017# => X"a65207ff",
		16#3018# => X"bc120000",
		16#3019# => X"0c0001c9",
		16#301a# => X"d4015830",
		16#301b# => X"8681006c",
		16#301c# => X"84410068",
		16#301d# => X"e0541000",
		16#301e# => X"9e420432",
		16#301f# => X"bdb20020",
		16#3020# => X"10000368",
		16#3021# => X"84810010",
		16#3022# => X"9d800040",
		16#3023# => X"9c420412",
		16#3024# => X"e18c9002",
		16#3025# => X"84610010",
		16#3026# => X"e19c6008",
		16#3027# => X"e0431048",
		16#3028# => X"e04c1004",
		16#3029# => X"a8620000",
		16#302a# => X"07ffecce",
		16#302b# => X"9e52fbcd",
		16#302c# => X"18c0fe10",
		16#302d# => X"aa0b0000",
		16#302e# => X"9ce00001",
		16#302f# => X"e2103000",
		16#3030# => X"a9cc0000",
		16#3031# => X"d4013858",
		16#3032# => X"a8500000",
		16#3033# => X"a86e0000",
		16#3034# => X"19800001",
		16#3035# => X"e0830004",
		16#3036# => X"e0620004",
		16#3037# => X"18400001",
		16#3038# => X"a98c4088",
		16#3039# => X"84ac0000",
		16#303a# => X"84cc0004",
		16#303b# => X"07ffe97c",
		16#303c# => X"a8424090",
		16#303d# => X"84a20000",
		16#303e# => X"84c20004",
		16#303f# => X"18400001",
		16#3040# => X"e06b0004",
		16#3041# => X"e08c0004",
		16#3042# => X"07ffe997",
		16#3043# => X"a8424098",
		16#3044# => X"84a20000",
		16#3045# => X"84c20004",
		16#3046# => X"e06b0004",
		16#3047# => X"e08c0004",
		16#3048# => X"07ffe950",
		16#3049# => X"18400001",
		16#304a# => X"a8720000",
		16#304b# => X"d4015808",
		16#304c# => X"d401600c",
		16#304d# => X"07ffec72",
		16#304e# => X"a84240a0",
		16#304f# => X"84a20000",
		16#3050# => X"84c20004",
		16#3051# => X"e06b0004",
		16#3052# => X"e08c0004",
		16#3053# => X"07ffe986",
		16#3054# => X"15000000",
		16#3055# => X"84610008",
		16#3056# => X"8481000c",
		16#3057# => X"e0ab0004",
		16#3058# => X"e0cc0004",
		16#3059# => X"07ffe93f",
		16#305a# => X"15000000",
		16#305b# => X"aa0b0000",
		16#305c# => X"a86c0000",
		16#305d# => X"a8500000",
		16#305e# => X"e0830004",
		16#305f# => X"e0620004",
		16#3060# => X"07ffece4",
		16#3061# => X"a9cc0000",
		16#3062# => X"18800001",
		16#3063# => X"a86e0000",
		16#3064# => X"a8844080",
		16#3065# => X"84a40000",
		16#3066# => X"84c40004",
		16#3067# => X"e0830004",
		16#3068# => X"e0620004",
		16#3069# => X"07ffebfe",
		16#306a# => X"d4015808",
		16#306b# => X"bd8b0000",
		16#306c# => X"0c000011",
		16#306d# => X"9ce00001",
		16#306e# => X"07ffec51",
		16#306f# => X"84610008",
		16#3070# => X"a9b00000",
		16#3071# => X"e06b0004",
		16#3072# => X"e08c0004",
		16#3073# => X"e0ad0004",
		16#3074# => X"e0ce0004",
		16#3075# => X"07ffeb98",
		16#3076# => X"15000000",
		16#3077# => X"bc2b0000",
		16#3078# => X"0c000005",
		16#3079# => X"9ce00001",
		16#307a# => X"84c10008",
		16#307b# => X"9cc6ffff",
		16#307c# => X"d4013008",
		16#307d# => X"84410008",
		16#307e# => X"bc420016",
		16#307f# => X"10000017",
		16#3080# => X"d401383c",
		16#3081# => X"18600001",
		16#3082# => X"b9c20003",
		16#3083# => X"85e10010",
		16#3084# => X"a8634118",
		16#3085# => X"a99c0000",
		16#3086# => X"a9af0000",
		16#3087# => X"e1ce1800",
		16#3088# => X"e0ac0004",
		16#3089# => X"e0cd0004",
		16#308a# => X"846e0000",
		16#308b# => X"848e0004",
		16#308c# => X"07ffeb9f",
		16#308d# => X"15000000",
		16#308e# => X"bd4b0000",
		16#308f# => X"0c0002fd",
		16#3090# => X"9ce00000",
		16#3091# => X"84810008",
		16#3092# => X"9cc00000",
		16#3093# => X"9c84ffff",
		16#3094# => X"d401303c",
		16#3095# => X"d4012008",
		16#3096# => X"9e94ffff",
		16#3097# => X"e2549002",
		16#3098# => X"bd720000",
		16#3099# => X"0c0002ea",
		16#309a# => X"9c600000",
		16#309b# => X"d4019024",
		16#309c# => X"d4011834",
		16#309d# => X"84810008",
		16#309e# => X"bd840000",
		16#309f# => X"100002db",
		16#30a0# => X"84c10024",
		16#30a1# => X"9ce00000",
		16#30a2# => X"e0c62000",
		16#30a3# => X"d4012048",
		16#30a4# => X"d4013024",
		16#30a5# => X"d4013840",
		16#30a6# => X"84e10000",
		16#30a7# => X"bc470009",
		16#30a8# => X"10000144",
		16#30a9# => X"9c400000",
		16#30aa# => X"bda70005",
		16#30ab# => X"10000005",
		16#30ac# => X"9dc00001",
		16#30ad# => X"9ce7fffc",
		16#30ae# => X"9dc00000",
		16#30af# => X"d4013800",
		16#30b0# => X"84410000",
		16#30b1# => X"bc020003",
		16#30b2# => X"100004bc",
		16#30b3# => X"bd420003",
		16#30b4# => X"0c0002e8",
		16#30b5# => X"bc020002",
		16#30b6# => X"84610000",
		16#30b7# => X"bc030004",
		16#30b8# => X"100004b9",
		16#30b9# => X"bc030005",
		16#30ba# => X"0c0002e4",
		16#30bb# => X"9cc0ffff",
		16#30bc# => X"9c800001",
		16#30bd# => X"d4012044",
		16#30be# => X"84c10008",
		16#30bf# => X"84e10018",
		16#30c0# => X"e0c63800",
		16#30c1# => X"9e260001",
		16#30c2# => X"bd510000",
		16#30c3# => X"0c0004e3",
		16#30c4# => X"d4013038",
		16#30c5# => X"d401881c",
		16#30c6# => X"9c400000",
		16#30c7# => X"bc510017",
		16#30c8# => X"0c00060b",
		16#30c9# => X"d41e1044",
		16#30ca# => X"9da00001",
		16#30cb# => X"9d800004",
		16#30cc# => X"e18c6000",
		16#30cd# => X"a84d0000",
		16#30ce# => X"9c6c0014",
		16#30cf# => X"e4a38800",
		16#30d0# => X"13fffffc",
		16#30d1# => X"9dad0001",
		16#30d2# => X"84c1001c",
		16#30d3# => X"d41e1044",
		16#30d4# => X"bca6000e",
		16#30d5# => X"10000003",
		16#30d6# => X"9d800001",
		16#30d7# => X"9d800000",
		16#30d8# => X"a87e0000",
		16#30d9# => X"a8820000",
		16#30da# => X"04000ccf",
		16#30db# => X"e1ce6003",
		16#30dc# => X"d4015820",
		16#30dd# => X"bc0e0000",
		16#30de# => X"0c00011f",
		16#30df# => X"d41e5840",
		16#30e0# => X"84c10008",
		16#30e1# => X"85a10068",
		16#30e2# => X"bda6000e",
		16#30e3# => X"10000003",
		16#30e4# => X"9d800001",
		16#30e5# => X"9d800000",
		16#30e6# => X"a58c00ff",
		16#30e7# => X"bc0c0000",
		16#30e8# => X"100001ee",
		16#30e9# => X"84410044",
		16#30ea# => X"bd8d0000",
		16#30eb# => X"100001ec",
		16#30ec# => X"bc020000",
		16#30ed# => X"84e10008",
		16#30ee# => X"18600001",
		16#30ef# => X"b9870003",
		16#30f0# => X"a8634118",
		16#30f1# => X"8441001c",
		16#30f2# => X"e18c1800",
		16#30f3# => X"bd420000",
		16#30f4# => X"84cc0000",
		16#30f5# => X"84ec0004",
		16#30f6# => X"d4013000",
		16#30f7# => X"d4013804",
		16#30f8# => X"10000007",
		16#30f9# => X"a9dc0000",
		16#30fa# => X"84e10018",
		16#30fb# => X"bd870000",
		16#30fc# => X"10000353",
		16#30fd# => X"84c1001c",
		16#30fe# => X"a9dc0000",
		16#30ff# => X"87810010",
		16#3100# => X"84410020",
		16#3101# => X"a8ee0000",
		16#3102# => X"a91c0000",
		16#3103# => X"9c420001",
		16#3104# => X"e0670004",
		16#3105# => X"e0880004",
		16#3106# => X"84a10000",
		16#3107# => X"84c10004",
		16#3108# => X"07ffe9d4",
		16#3109# => X"d4011028",
		16#310a# => X"e06b0004",
		16#310b# => X"e08c0004",
		16#310c# => X"07ffec38",
		16#310d# => X"15000000",
		16#310e# => X"a86b0000",
		16#310f# => X"07ffebb0",
		16#3110# => X"aa4b0000",
		16#3111# => X"84a10000",
		16#3112# => X"84c10004",
		16#3113# => X"e06b0004",
		16#3114# => X"e08c0004",
		16#3115# => X"07ffe8c4",
		16#3116# => X"15000000",
		16#3117# => X"a8ee0000",
		16#3118# => X"a91c0000",
		16#3119# => X"e0ab0004",
		16#311a# => X"e0cc0004",
		16#311b# => X"e0670004",
		16#311c# => X"e0880004",
		16#311d# => X"07ffe89a",
		16#311e# => X"15000000",
		16#311f# => X"84610020",
		16#3120# => X"a9ac0000",
		16#3121# => X"9d920030",
		16#3122# => X"a9cb0000",
		16#3123# => X"d8036000",
		16#3124# => X"a8ee0000",
		16#3125# => X"8481001c",
		16#3126# => X"bc040001",
		16#3127# => X"1000005c",
		16#3128# => X"a98d0000",
		16#3129# => X"1b000001",
		16#312a# => X"a8ee0000",
		16#312b# => X"a90d0000",
		16#312c# => X"ab1840b0",
		16#312d# => X"e0670004",
		16#312e# => X"e0880004",
		16#312f# => X"84b80000",
		16#3130# => X"84d80004",
		16#3131# => X"07ffe8a8",
		16#3132# => X"18400001",
		16#3133# => X"a9cb0000",
		16#3134# => X"a90c0000",
		16#3135# => X"a8ee0000",
		16#3136# => X"a8424080",
		16#3137# => X"aa0c0000",
		16#3138# => X"84a20000",
		16#3139# => X"84c20004",
		16#313a# => X"e0670004",
		16#313b# => X"e0880004",
		16#313c# => X"07ffead1",
		16#313d# => X"9e400001",
		16#313e# => X"bc2b0000",
		16#313f# => X"10000004",
		16#3140# => X"a65200ff",
		16#3141# => X"aa4b0000",
		16#3142# => X"a65200ff",
		16#3143# => X"bc120000",
		16#3144# => X"10000182",
		16#3145# => X"9e800001",
		16#3146# => X"8781001c",
		16#3147# => X"00000017",
		16#3148# => X"86c10028",
		16#3149# => X"84b80000",
		16#314a# => X"84d80004",
		16#314b# => X"07ffe88e",
		16#314c# => X"15000000",
		16#314d# => X"18e00001",
		16#314e# => X"a9cb0000",
		16#314f# => X"a8e74080",
		16#3150# => X"a86e0000",
		16#3151# => X"a88c0000",
		16#3152# => X"84a70000",
		16#3153# => X"84c70004",
		16#3154# => X"07ffeab9",
		16#3155# => X"aa0c0000",
		16#3156# => X"bc2b0000",
		16#3157# => X"10000004",
		16#3158# => X"a75a00ff",
		16#3159# => X"ab4b0000",
		16#315a# => X"a75a00ff",
		16#315b# => X"bc1a0000",
		16#315c# => X"100004ce",
		16#315d# => X"15000000",
		16#315e# => X"a86e0000",
		16#315f# => X"84a10000",
		16#3160# => X"84c10004",
		16#3161# => X"07ffe97b",
		16#3162# => X"a8900000",
		16#3163# => X"e06b0004",
		16#3164# => X"e08c0004",
		16#3165# => X"07ffebdf",
		16#3166# => X"a84e0000",
		16#3167# => X"a86b0000",
		16#3168# => X"07ffeb57",
		16#3169# => X"aa4b0000",
		16#316a# => X"84a10000",
		16#316b# => X"84c10004",
		16#316c# => X"e06b0004",
		16#316d# => X"e08c0004",
		16#316e# => X"07ffe86b",
		16#316f# => X"9e940001",
		16#3170# => X"a8700000",
		16#3171# => X"e0ab0004",
		16#3172# => X"e0cc0004",
		16#3173# => X"e0830004",
		16#3174# => X"e0620004",
		16#3175# => X"07ffe842",
		16#3176# => X"9f400001",
		16#3177# => X"a88b0000",
		16#3178# => X"a8440000",
		16#3179# => X"9c920030",
		16#317a# => X"a86c0000",
		16#317b# => X"d8162000",
		16#317c# => X"e0830004",
		16#317d# => X"e0620004",
		16#317e# => X"e41ca000",
		16#317f# => X"0fffffca",
		16#3180# => X"9ed60001",
		16#3181# => X"d401b028",
		16#3182# => X"a8eb0000",
		16#3183# => X"a9a70000",
		16#3184# => X"a9cc0000",
		16#3185# => X"a8c70000",
		16#3186# => X"a8ec0000",
		16#3187# => X"e06d0004",
		16#3188# => X"e08e0004",
		16#3189# => X"e0a60004",
		16#318a# => X"e0c70004",
		16#318b# => X"07ffe80d",
		16#318c# => X"15000000",
		16#318d# => X"aa0b0000",
		16#318e# => X"a8ec0000",
		16#318f# => X"a8d00000",
		16#3190# => X"84410008",
		16#3191# => X"a9cc0000",
		16#3192# => X"84610000",
		16#3193# => X"84810004",
		16#3194# => X"e0a60004",
		16#3195# => X"e0c70004",
		16#3196# => X"07ffead1",
		16#3197# => X"d401105c",
		16#3198# => X"bd8b0000",
		16#3199# => X"10000013",
		16#319a# => X"84610028",
		16#319b# => X"a8ee0000",
		16#319c# => X"a8d00000",
		16#319d# => X"84610000",
		16#319e# => X"84810004",
		16#319f# => X"e0a60004",
		16#31a0# => X"e0c70004",
		16#31a1# => X"07ffea4e",
		16#31a2# => X"15000000",
		16#31a3# => X"bc0b0000",
		16#31a4# => X"0c000123",
		16#31a5# => X"a87e0000",
		16#31a6# => X"84610008",
		16#31a7# => X"a6520001",
		16#31a8# => X"bc320000",
		16#31a9# => X"0c00011d",
		16#31aa# => X"d401185c",
		16#31ab# => X"84610028",
		16#31ac# => X"00000003",
		16#31ad# => X"84810020",
		16#31ae# => X"a8620000",
		16#31af# => X"9c43ffff",
		16#31b0# => X"90c20000",
		16#31b1# => X"bc060039",
		16#31b2# => X"0c000498",
		16#31b3# => X"e4222000",
		16#31b4# => X"13fffffa",
		16#31b5# => X"9ce00030",
		16#31b6# => X"d4012020",
		16#31b7# => X"8481005c",
		16#31b8# => X"84c10020",
		16#31b9# => X"9c840001",
		16#31ba# => X"d4011828",
		16#31bb# => X"d4012008",
		16#31bc# => X"d8063800",
		16#31bd# => X"9cc00031",
		16#31be# => X"00000108",
		16#31bf# => X"d8023000",
		16#31c0# => X"9c40270f",
		16#31c1# => X"84e10014",
		16#31c2# => X"19600001",
		16#31c3# => X"d4071000",
		16#31c4# => X"84410010",
		16#31c5# => X"bc220000",
		16#31c6# => X"1000000b",
		16#31c7# => X"a96b4079",
		16#31c8# => X"1860000f",
		16#31c9# => X"19600001",
		16#31ca# => X"a863ffff",
		16#31cb# => X"e09c1803",
		16#31cc# => X"bc040000",
		16#31cd# => X"10000004",
		16#31ce# => X"a96b4070",
		16#31cf# => X"19600001",
		16#31d0# => X"a96b4079",
		16#31d1# => X"848100a0",
		16#31d2# => X"bc040000",
		16#31d3# => X"13fffe29",
		16#31d4# => X"9c4b0003",
		16#31d5# => X"90620000",
		16#31d6# => X"bc030000",
		16#31d7# => X"10000003",
		16#31d8# => X"84c100a0",
		16#31d9# => X"9c4b0008",
		16#31da# => X"03fffe22",
		16#31db# => X"d4061000",
		16#31dc# => X"18607fff",
		16#31dd# => X"9c400001",
		16#31de# => X"a863ffff",
		16#31df# => X"d40e1000",
		16#31e0# => X"03fffdfb",
		16#31e1# => X"e39c1803",
		16#31e2# => X"18c0000f",
		16#31e3# => X"18e03ff0",
		16#31e4# => X"a8c6ffff",
		16#31e5# => X"9c400000",
		16#31e6# => X"e2103003",
		16#31e7# => X"9e52fc01",
		16#31e8# => X"e2103804",
		16#31e9# => X"8681006c",
		16#31ea# => X"03fffe48",
		16#31eb# => X"d4011058",
		16#31ec# => X"9c60ffff",
		16#31ed# => X"9c800001",
		16#31ee# => X"d4011000",
		16#31ef# => X"d4011838",
		16#31f0# => X"a9c20000",
		16#31f1# => X"d4012044",
		16#31f2# => X"d401181c",
		16#31f3# => X"d4011018",
		16#31f4# => X"9c400000",
		16#31f5# => X"d41e1044",
		16#31f6# => X"a87e0000",
		16#31f7# => X"04000bb2",
		16#31f8# => X"a8820000",
		16#31f9# => X"d4015820",
		16#31fa# => X"bc0e0000",
		16#31fb# => X"13fffee5",
		16#31fc# => X"d41e5840",
		16#31fd# => X"84e10010",
		16#31fe# => X"84410008",
		16#31ff# => X"d401382c",
		16#3200# => X"bda20000",
		16#3201# => X"100002b6",
		16#3202# => X"aa5c0000",
		16#3203# => X"a5e2000f",
		16#3204# => X"18600001",
		16#3205# => X"ba020084",
		16#3206# => X"b9ef0003",
		16#3207# => X"a8634118",
		16#3208# => X"a5d00010",
		16#3209# => X"e1af1800",
		16#320a# => X"9f400002",
		16#320b# => X"bc0e0000",
		16#320c# => X"86cd0000",
		16#320d# => X"0c000181",
		16#320e# => X"868d0004",
		16#320f# => X"bc100000",
		16#3210# => X"10000014",
		16#3211# => X"a9760000",
		16#3212# => X"1b000001",
		16#3213# => X"ab1841e0",
		16#3214# => X"a9940000",
		16#3215# => X"a4500001",
		16#3216# => X"a86b0000",
		16#3217# => X"a88c0000",
		16#3218# => X"bc020000",
		16#3219# => X"10000006",
		16#321a# => X"ba100081",
		16#321b# => X"84b80000",
		16#321c# => X"84d80004",
		16#321d# => X"07ffe7bc",
		16#321e# => X"9f5a0001",
		16#321f# => X"bc300000",
		16#3220# => X"13fffff5",
		16#3221# => X"9f180008",
		16#3222# => X"aacb0000",
		16#3223# => X"aa8c0000",
		16#3224# => X"8581002c",
		16#3225# => X"a8520000",
		16#3226# => X"a9b60000",
		16#3227# => X"a86c0000",
		16#3228# => X"a9d40000",
		16#3229# => X"e0830004",
		16#322a# => X"e0620004",
		16#322b# => X"e0ad0004",
		16#322c# => X"e0ce0004",
		16#322d# => X"07ffe8af",
		16#322e# => X"15000000",
		16#322f# => X"aa4b0000",
		16#3230# => X"d401602c",
		16#3231# => X"84e1003c",
		16#3232# => X"bc070000",
		16#3233# => X"1000003c",
		16#3234# => X"a8520000",
		16#3235# => X"85c1002c",
		16#3236# => X"a86e0000",
		16#3237# => X"19c00001",
		16#3238# => X"e0830004",
		16#3239# => X"e0620004",
		16#323a# => X"a9ce40a8",
		16#323b# => X"84ae0000",
		16#323c# => X"84ce0004",
		16#323d# => X"07ffea2a",
		16#323e# => X"15000000",
		16#323f# => X"bd6b0000",
		16#3240# => X"1000002f",
		16#3241# => X"8441001c",
		16#3242# => X"bda20000",
		16#3243# => X"1000002c",
		16#3244# => X"84610038",
		16#3245# => X"bda30000",
		16#3246# => X"13fffe9a",
		16#3247# => X"8581002c",
		16#3248# => X"1b000001",
		16#3249# => X"a9b20000",
		16#324a# => X"a9cc0000",
		16#324b# => X"ab1840b0",
		16#324c# => X"e06d0004",
		16#324d# => X"e08e0004",
		16#324e# => X"84b80000",
		16#324f# => X"84d80004",
		16#3250# => X"07ffe789",
		16#3251# => X"1840fcc0",
		16#3252# => X"84810008",
		16#3253# => X"9c7a0001",
		16#3254# => X"9c84ffff",
		16#3255# => X"aa4b0000",
		16#3256# => X"d401205c",
		16#3257# => X"07ffea68",
		16#3258# => X"d401602c",
		16#3259# => X"85a1002c",
		16#325a# => X"84e10038",
		16#325b# => X"a9ed0000",
		16#325c# => X"a9d20000",
		16#325d# => X"e0ab0004",
		16#325e# => X"e0cc0004",
		16#325f# => X"e06e0004",
		16#3260# => X"e08f0004",
		16#3261# => X"07ffe778",
		16#3262# => X"d401384c",
		16#3263# => X"1a600001",
		16#3264# => X"e06b0004",
		16#3265# => X"e08c0004",
		16#3266# => X"aa7340b8",
		16#3267# => X"84b30000",
		16#3268# => X"84d30004",
		16#3269# => X"07ffe72f",
		16#326a# => X"15000000",
		16#326b# => X"aa8b0000",
		16#326c# => X"a9cc0000",
		16#326d# => X"00000140",
		16#326e# => X"e3541000",
		16#326f# => X"07ffea50",
		16#3270# => X"a87a0000",
		16#3271# => X"85e1002c",
		16#3272# => X"a9b20000",
		16#3273# => X"a9cf0000",
		16#3274# => X"e06b0004",
		16#3275# => X"e08c0004",
		16#3276# => X"e0ad0004",
		16#3277# => X"e0ce0004",
		16#3278# => X"07ffe761",
		16#3279# => X"15000000",
		16#327a# => X"19a00001",
		16#327b# => X"e06b0004",
		16#327c# => X"e08c0004",
		16#327d# => X"a9ad40b8",
		16#327e# => X"84ad0000",
		16#327f# => X"84cd0004",
		16#3280# => X"07ffe718",
		16#3281# => X"15000000",
		16#3282# => X"1860fcc0",
		16#3283# => X"a9ab0000",
		16#3284# => X"8481001c",
		16#3285# => X"ab0c0000",
		16#3286# => X"e34d1800",
		16#3287# => X"bc240000",
		16#3288# => X"10000121",
		16#3289# => X"a9cc0000",
		16#328a# => X"85e1002c",
		16#328b# => X"a8520000",
		16#328c# => X"a86f0000",
		16#328d# => X"19e00001",
		16#328e# => X"e0830004",
		16#328f# => X"e0620004",
		16#3290# => X"a9ef40c0",
		16#3291# => X"84af0000",
		16#3292# => X"84cf0004",
		16#3293# => X"07ffe724",
		16#3294# => X"aa180000",
		16#3295# => X"aacb0000",
		16#3296# => X"a9fa0000",
		16#3297# => X"aa760000",
		16#3298# => X"aa8c0000",
		16#3299# => X"e0730004",
		16#329a# => X"e0940004",
		16#329b# => X"e0af0004",
		16#329c# => X"e0d00004",
		16#329d# => X"07ffe98e",
		16#329e# => X"a9cc0000",
		16#329f# => X"bd4b0000",
		16#32a0# => X"100001c5",
		16#32a1# => X"18c08000",
		16#32a2# => X"a9f60000",
		16#32a3# => X"e2ba3000",
		16#32a4# => X"aa0e0000",
		16#32a5# => X"a9b50000",
		16#32a6# => X"a9d80000",
		16#32a7# => X"e06f0004",
		16#32a8# => X"e0900004",
		16#32a9# => X"e0ad0004",
		16#32aa# => X"e0ce0004",
		16#32ab# => X"07ffe9bc",
		16#32ac# => X"15000000",
		16#32ad# => X"bd8b0000",
		16#32ae# => X"0ffffe33",
		16#32af# => X"84c10008",
		16#32b0# => X"8441001c",
		16#32b1# => X"aa420000",
		16#32b2# => X"84810018",
		16#32b3# => X"84c10020",
		16#32b4# => X"ac84ffff",
		16#32b5# => X"d4013028",
		16#32b6# => X"d4012008",
		16#32b7# => X"9dc00000",
		16#32b8# => X"a87e0000",
		16#32b9# => X"04000b1d",
		16#32ba# => X"a8820000",
		16#32bb# => X"bc120000",
		16#32bc# => X"1000000a",
		16#32bd# => X"e0ce9005",
		16#32be# => X"e0e03002",
		16#32bf# => X"e0c73004",
		16#32c0# => X"bd660000",
		16#32c1# => X"0c0001e2",
		16#32c2# => X"e0c07002",
		16#32c3# => X"a87e0000",
		16#32c4# => X"04000b12",
		16#32c5# => X"a8920000",
		16#32c6# => X"a87e0000",
		16#32c7# => X"04000b0f",
		16#32c8# => X"84810030",
		16#32c9# => X"84610028",
		16#32ca# => X"9c800000",
		16#32cb# => X"84e10008",
		16#32cc# => X"d8032000",
		16#32cd# => X"9c470001",
		16#32ce# => X"84c10014",
		16#32cf# => X"84e100a0",
		16#32d0# => X"d4061000",
		16#32d1# => X"bc070000",
		16#32d2# => X"13fffd2a",
		16#32d3# => X"85610020",
		16#32d4# => X"03fffd28",
		16#32d5# => X"d4071800",
		16#32d6# => X"bc020000",
		16#32d7# => X"100000ce",
		16#32d8# => X"84610000",
		16#32d9# => X"bd430001",
		16#32da# => X"0c000368",
		16#32db# => X"84c1001c",
		16#32dc# => X"84e10040",
		16#32dd# => X"9e06ffff",
		16#32de# => X"e5878000",
		16#32df# => X"10000353",
		16#32e0# => X"84410040",
		16#32e1# => X"e2078002",
		16#32e2# => X"8481001c",
		16#32e3# => X"bd640000",
		16#32e4# => X"0c000375",
		16#32e5# => X"84c10034",
		16#32e6# => X"85c10034",
		16#32e7# => X"85a1001c",
		16#32e8# => X"84e10034",
		16#32e9# => X"84410024",
		16#32ea# => X"e0e76800",
		16#32eb# => X"e0426800",
		16#32ec# => X"a87e0000",
		16#32ed# => X"9c800001",
		16#32ee# => X"d4013834",
		16#32ef# => X"04000be7",
		16#32f0# => X"d4011024",
		16#32f1# => X"aa4b0000",
		16#32f2# => X"84610024",
		16#32f3# => X"bda30000",
		16#32f4# => X"1000000f",
		16#32f5# => X"bdae0000",
		16#32f6# => X"1000000e",
		16#32f7# => X"84e10040",
		16#32f8# => X"e5a37000",
		16#32f9# => X"10000003",
		16#32fa# => X"a9830000",
		16#32fb# => X"a98e0000",
		16#32fc# => X"84810034",
		16#32fd# => X"84c10024",
		16#32fe# => X"e0846002",
		16#32ff# => X"e0c66002",
		16#3300# => X"d4012034",
		16#3301# => X"e1ce6002",
		16#3302# => X"d4013024",
		16#3303# => X"84e10040",
		16#3304# => X"bda70000",
		16#3305# => X"10000018",
		16#3306# => X"84410044",
		16#3307# => X"bc020000",
		16#3308# => X"10000324",
		16#3309# => X"bdb00000",
		16#330a# => X"1000000e",
		16#330b# => X"a8920000",
		16#330c# => X"a87e0000",
		16#330d# => X"04000c67",
		16#330e# => X"a8b00000",
		16#330f# => X"a87e0000",
		16#3310# => X"a88b0000",
		16#3311# => X"84a10030",
		16#3312# => X"04000bd1",
		16#3313# => X"aa4b0000",
		16#3314# => X"84810030",
		16#3315# => X"a87e0000",
		16#3316# => X"04000ac0",
		16#3317# => X"d4015830",
		16#3318# => X"84610040",
		16#3319# => X"e2038002",
		16#331a# => X"bc100000",
		16#331b# => X"0c00031f",
		16#331c# => X"a87e0000",
		16#331d# => X"9c800001",
		16#331e# => X"04000bb8",
		16#331f# => X"a87e0000",
		16#3320# => X"84810048",
		16#3321# => X"bda40000",
		16#3322# => X"10000007",
		16#3323# => X"a84b0000",
		16#3324# => X"a87e0000",
		16#3325# => X"a88b0000",
		16#3326# => X"04000c4e",
		16#3327# => X"84a10048",
		16#3328# => X"a84b0000",
		16#3329# => X"84c10000",
		16#332a# => X"bd460001",
		16#332b# => X"0c000282",
		16#332c# => X"9e000000",
		16#332d# => X"84610048",
		16#332e# => X"bc030000",
		16#332f# => X"0c000269",
		16#3330# => X"9da00001",
		16#3331# => X"84810024",
		16#3332# => X"e1ad2000",
		16#3333# => X"a5ad001f",
		16#3334# => X"bc0d0000",
		16#3335# => X"0c000176",
		16#3336# => X"9d80001c",
		16#3337# => X"84e10034",
		16#3338# => X"84610024",
		16#3339# => X"e0e76000",
		16#333a# => X"e0636000",
		16#333b# => X"d4013834",
		16#333c# => X"e1ce6000",
		16#333d# => X"d4011824",
		16#333e# => X"84810034",
		16#333f# => X"bda40000",
		16#3340# => X"10000008",
		16#3341# => X"84c10024",
		16#3342# => X"a87e0000",
		16#3343# => X"84810030",
		16#3344# => X"04000c88",
		16#3345# => X"84a10034",
		16#3346# => X"d4015830",
		16#3347# => X"84c10024",
		16#3348# => X"bda60000",
		16#3349# => X"10000008",
		16#334a# => X"84e1003c",
		16#334b# => X"a8820000",
		16#334c# => X"a87e0000",
		16#334d# => X"04000c7f",
		16#334e# => X"a8a60000",
		16#334f# => X"a84b0000",
		16#3350# => X"84e1003c",
		16#3351# => X"bc070000",
		16#3352# => X"0c00022b",
		16#3353# => X"15000000",
		16#3354# => X"84c1001c",
		16#3355# => X"bd460000",
		16#3356# => X"10000112",
		16#3357# => X"84e10044",
		16#3358# => X"84e10000",
		16#3359# => X"bd470002",
		16#335a# => X"10000003",
		16#335b# => X"9d800001",
		16#335c# => X"9d800000",
		16#335d# => X"a58c00ff",
		16#335e# => X"bc0c0000",
		16#335f# => X"10000109",
		16#3360# => X"84e10044",
		16#3361# => X"8461001c",
		16#3362# => X"bc230000",
		16#3363# => X"13ffff4f",
		16#3364# => X"a8c30000",
		16#3365# => X"a8820000",
		16#3366# => X"9ca00005",
		16#3367# => X"04000a7b",
		16#3368# => X"a87e0000",
		16#3369# => X"84610030",
		16#336a# => X"a88b0000",
		16#336b# => X"04000cc0",
		16#336c# => X"a84b0000",
		16#336d# => X"bd4b0000",
		16#336e# => X"0fffff44",
		16#336f# => X"15000000",
		16#3370# => X"84e10020",
		16#3371# => X"9c600031",
		16#3372# => X"9c870001",
		16#3373# => X"d8071800",
		16#3374# => X"d4012028",
		16#3375# => X"84c10008",
		16#3376# => X"9dc00000",
		16#3377# => X"9cc60001",
		16#3378# => X"03ffff40",
		16#3379# => X"d4013008",
		16#337a# => X"84410034",
		16#337b# => X"84610008",
		16#337c# => X"9cc00000",
		16#337d# => X"e0421802",
		16#337e# => X"e0801802",
		16#337f# => X"d4011034",
		16#3380# => X"d4012040",
		16#3381# => X"03fffd25",
		16#3382# => X"d4013048",
		16#3383# => X"e2409002",
		16#3384# => X"9c400000",
		16#3385# => X"d4019034",
		16#3386# => X"03fffd17",
		16#3387# => X"d4011024",
		16#3388# => X"9c400020",
		16#3389# => X"e0429002",
		16#338a# => X"03fffc9f",
		16#338b# => X"e0441008",
		16#338c# => X"03fffd0a",
		16#338d# => X"d401383c",
		16#338e# => X"19800001",
		16#338f# => X"a8670000",
		16#3390# => X"a98c41e0",
		16#3391# => X"a85c0000",
		16#3392# => X"84ac0020",
		16#3393# => X"84cc0024",
		16#3394# => X"e0830004",
		16#3395# => X"e0620004",
		16#3396# => X"07ffe746",
		16#3397# => X"a610000f",
		16#3398# => X"9f400003",
		16#3399# => X"aa4b0000",
		16#339a# => X"03fffe75",
		16#339b# => X"d401602c",
		16#339c# => X"100001de",
		16#339d# => X"9cc0ffff",
		16#339e# => X"9dc00000",
		16#339f# => X"9ce00001",
		16#33a0# => X"d4013038",
		16#33a1# => X"d4013844",
		16#33a2# => X"d401301c",
		16#33a3# => X"03fffe51",
		16#33a4# => X"d4017018",
		16#33a5# => X"86010040",
		16#33a6# => X"85c10034",
		16#33a7# => X"03ffff4b",
		16#33a8# => X"86410044",
		16#33a9# => X"84e10008",
		16#33aa# => X"8441001c",
		16#33ab# => X"d401385c",
		16#33ac# => X"d401104c",
		16#33ad# => X"84610044",
		16#33ae# => X"bc030000",
		16#33af# => X"10000136",
		16#33b0# => X"8481004c",
		16#33b1# => X"18c00001",
		16#33b2# => X"9e64ffff",
		16#33b3# => X"a8c64118",
		16#33b4# => X"ba730003",
		16#33b5# => X"e1933000",
		16#33b6# => X"1a600001",
		16#33b7# => X"84ac0000",
		16#33b8# => X"84cc0004",
		16#33b9# => X"aa7340c8",
		16#33ba# => X"84730000",
		16#33bb# => X"84930004",
		16#33bc# => X"07ffe720",
		16#33bd# => X"aada0000",
		16#33be# => X"84e10020",
		16#33bf# => X"aaee0000",
		16#33c0# => X"9ce70001",
		16#33c1# => X"e0b60004",
		16#33c2# => X"e0d70004",
		16#33c3# => X"e06b0004",
		16#33c4# => X"e08c0004",
		16#33c5# => X"07ffe5f2",
		16#33c6# => X"d4013828",
		16#33c7# => X"8461002c",
		16#33c8# => X"aab20000",
		16#33c9# => X"aac30000",
		16#33ca# => X"aa0c0000",
		16#33cb# => X"e0750004",
		16#33cc# => X"e0960004",
		16#33cd# => X"07ffe977",
		16#33ce# => X"aa8b0000",
		16#33cf# => X"a86b0000",
		16#33d0# => X"07ffe8ef",
		16#33d1# => X"a84b0000",
		16#33d2# => X"85e1002c",
		16#33d3# => X"aab20000",
		16#33d4# => X"aacf0000",
		16#33d5# => X"e0ab0004",
		16#33d6# => X"e0cc0004",
		16#33d7# => X"e0750004",
		16#33d8# => X"e0960004",
		16#33d9# => X"07ffe5de",
		16#33da# => X"aad00000",
		16#33db# => X"9ce20030",
		16#33dc# => X"ab4b0000",
		16#33dd# => X"84410020",
		16#33de# => X"aab40000",
		16#33df# => X"a9ba0000",
		16#33e0# => X"a9cc0000",
		16#33e1# => X"d8023800",
		16#33e2# => X"e0750004",
		16#33e3# => X"e0960004",
		16#33e4# => X"e0ad0004",
		16#33e5# => X"e0ce0004",
		16#33e6# => X"07ffe845",
		16#33e7# => X"aa4c0000",
		16#33e8# => X"bd4b0000",
		16#33e9# => X"100002e7",
		16#33ea# => X"18c00001",
		16#33eb# => X"a9ba0000",
		16#33ec# => X"a8c640a8",
		16#33ed# => X"84660000",
		16#33ee# => X"84860004",
		16#33ef# => X"e0ad0004",
		16#33f0# => X"e0ce0004",
		16#33f1# => X"07ffe5c6",
		16#33f2# => X"a9d00000",
		16#33f3# => X"a9b40000",
		16#33f4# => X"e0ab0004",
		16#33f5# => X"e0cc0004",
		16#33f6# => X"e06d0004",
		16#33f7# => X"e08e0004",
		16#33f8# => X"07ffe833",
		16#33f9# => X"15000000",
		16#33fa# => X"bd4b0000",
		16#33fb# => X"13fffdb0",
		16#33fc# => X"84e1004c",
		16#33fd# => X"bda70001",
		16#33fe# => X"13fffce2",
		16#33ff# => X"1b000001",
		16#3400# => X"9ec00001",
		16#3401# => X"ab1840b0",
		16#3402# => X"d401f060",
		16#3403# => X"85d80000",
		16#3404# => X"87180004",
		16#3405# => X"d401e064",
		16#3406# => X"d401c050",
		16#3407# => X"ab960000",
		16#3408# => X"d401c054",
		16#3409# => X"d401702c",
		16#340a# => X"aad00000",
		16#340b# => X"abce0000",
		16#340c# => X"00000014",
		16#340d# => X"87010028",
		16#340e# => X"18400001",
		16#340f# => X"a84240a8",
		16#3410# => X"84620000",
		16#3411# => X"84820004",
		16#3412# => X"07ffe5a5",
		16#3413# => X"15000000",
		16#3414# => X"a8b40000",
		16#3415# => X"e06b0004",
		16#3416# => X"e08c0004",
		16#3417# => X"07ffe850",
		16#3418# => X"a8d60000",
		16#3419# => X"bd8b0000",
		16#341a# => X"10000239",
		16#341b# => X"a8780000",
		16#341c# => X"8461004c",
		16#341d# => X"e57c1800",
		16#341e# => X"10000238",
		16#341f# => X"15000000",
		16#3420# => X"a8740000",
		16#3421# => X"a8960000",
		16#3422# => X"84c10054",
		16#3423# => X"a8be0000",
		16#3424# => X"07ffe5b5",
		16#3425# => X"9f9c0001",
		16#3426# => X"84a1002c",
		16#3427# => X"84c10050",
		16#3428# => X"a87a0000",
		16#3429# => X"a8920000",
		16#342a# => X"aa8b0000",
		16#342b# => X"07ffe5ae",
		16#342c# => X"aacc0000",
		16#342d# => X"aa4b0000",
		16#342e# => X"a88c0000",
		16#342f# => X"a8720000",
		16#3430# => X"07ffe914",
		16#3431# => X"aa0c0000",
		16#3432# => X"a86b0000",
		16#3433# => X"07ffe88c",
		16#3434# => X"a9cb0000",
		16#3435# => X"a8520000",
		16#3436# => X"a8700000",
		16#3437# => X"e0ab0004",
		16#3438# => X"e0cc0004",
		16#3439# => X"e0830004",
		16#343a# => X"e0620004",
		16#343b# => X"07ffe57c",
		16#343c# => X"9dce0030",
		16#343d# => X"ab4b0000",
		16#343e# => X"a8b40000",
		16#343f# => X"d8187000",
		16#3440# => X"a8d60000",
		16#3441# => X"a87a0000",
		16#3442# => X"a88c0000",
		16#3443# => X"07ffe824",
		16#3444# => X"aa4c0000",
		16#3445# => X"9f180001",
		16#3446# => X"a8ba0000",
		16#3447# => X"bd8b0000",
		16#3448# => X"0fffffc6",
		16#3449# => X"a8d20000",
		16#344a# => X"84c1005c",
		16#344b# => X"d401c028",
		16#344c# => X"87c10060",
		16#344d# => X"03fffe79",
		16#344e# => X"d4013008",
		16#344f# => X"bc260000",
		16#3450# => X"100001ef",
		16#3451# => X"19800001",
		16#3452# => X"84610000",
		16#3453# => X"84810004",
		16#3454# => X"a98c40c0",
		16#3455# => X"84ac0000",
		16#3456# => X"84cc0004",
		16#3457# => X"07ffe582",
		16#3458# => X"a9dc0000",
		16#3459# => X"87810010",
		16#345a# => X"e06b0004",
		16#345b# => X"e08c0004",
		16#345c# => X"a9bc0000",
		16#345d# => X"a98e0000",
		16#345e# => X"e0ac0004",
		16#345f# => X"e0cd0004",
		16#3460# => X"07ffe7e9",
		16#3461# => X"15000000",
		16#3462# => X"bd6b0000",
		16#3463# => X"13fffe4d",
		16#3464# => X"15000000",
		16#3465# => X"8441001c",
		16#3466# => X"03ffff0a",
		16#3467# => X"aa420000",
		16#3468# => X"bc270000",
		16#3469# => X"1000015b",
		16#346a# => X"bdae0000",
		16#346b# => X"84610020",
		16#346c# => X"9dc00001",
		16#346d# => X"d4011828",
		16#346e# => X"8601001c",
		16#346f# => X"86c10030",
		16#3470# => X"00000005",
		16#3471# => X"aa830000",
		16#3472# => X"04000970",
		16#3473# => X"9dce0001",
		16#3474# => X"aacb0000",
		16#3475# => X"a8760000",
		16#3476# => X"07fffaa8",
		16#3477# => X"a8820000",
		16#3478# => X"9d6b0030",
		16#3479# => X"a87e0000",
		16#347a# => X"d8145800",
		16#347b# => X"a8960000",
		16#347c# => X"9ca0000a",
		16#347d# => X"9cc00000",
		16#347e# => X"e56e8000",
		16#347f# => X"0ffffff3",
		16#3480# => X"9e940001",
		16#3481# => X"aa0b0000",
		16#3482# => X"d401b030",
		16#3483# => X"d401a028",
		16#3484# => X"9dc00000",
		16#3485# => X"9ca00001",
		16#3486# => X"a87e0000",
		16#3487# => X"04000b45",
		16#3488# => X"84810030",
		16#3489# => X"a8820000",
		16#348a# => X"a86b0000",
		16#348b# => X"04000ba0",
		16#348c# => X"d4015830",
		16#348d# => X"bd4b0000",
		16#348e# => X"0c0001e6",
		16#348f# => X"bc2b0000",
		16#3490# => X"84610028",
		16#3491# => X"00000003",
		16#3492# => X"84810020",
		16#3493# => X"a8660000",
		16#3494# => X"9cc3ffff",
		16#3495# => X"90e60000",
		16#3496# => X"bc070039",
		16#3497# => X"0c0001ed",
		16#3498# => X"e4262000",
		16#3499# => X"13fffffa",
		16#349a# => X"15000000",
		16#349b# => X"84c10008",
		16#349c# => X"d4011828",
		16#349d# => X"9cc60001",
		16#349e# => X"9c600031",
		16#349f# => X"84e10020",
		16#34a0# => X"d4013008",
		16#34a1# => X"03fffe17",
		16#34a2# => X"d8071800",
		16#34a3# => X"e0ce3004",
		16#34a4# => X"bd660000",
		16#34a5# => X"13fffe1e",
		16#34a6# => X"a87e0000",
		16#34a7# => X"0400092f",
		16#34a8# => X"a88e0000",
		16#34a9# => X"03fffe1b",
		16#34aa# => X"a87e0000",
		16#34ab# => X"9d800020",
		16#34ac# => X"e18c6802",
		16#34ad# => X"bdac0004",
		16#34ae# => X"1000022d",
		16#34af# => X"84c10034",
		16#34b0# => X"9d8cfffc",
		16#34b1# => X"e0846000",
		16#34b2# => X"e0c66000",
		16#34b3# => X"e1ce6000",
		16#34b4# => X"d4013034",
		16#34b5# => X"03fffe89",
		16#34b6# => X"d4012024",
		16#34b7# => X"84810008",
		16#34b8# => X"e2002002",
		16#34b9# => X"bc100000",
		16#34ba# => X"13fffd77",
		16#34bb# => X"9f400002",
		16#34bc# => X"a5f0000f",
		16#34bd# => X"18c00001",
		16#34be# => X"b9ef0003",
		16#34bf# => X"86610010",
		16#34c0# => X"a8c64118",
		16#34c1# => X"a99c0000",
		16#34c2# => X"e1ef3000",
		16#34c3# => X"a9b30000",
		16#34c4# => X"e06c0004",
		16#34c5# => X"e08d0004",
		16#34c6# => X"84af0000",
		16#34c7# => X"84cf0004",
		16#34c8# => X"07ffe511",
		16#34c9# => X"ba100084",
		16#34ca# => X"d401602c",
		16#34cb# => X"bc100000",
		16#34cc# => X"13fffd65",
		16#34cd# => X"aa4b0000",
		16#34ce# => X"1a800001",
		16#34cf# => X"a9d20000",
		16#34d0# => X"aa9441e0",
		16#34d1# => X"a9ac0000",
		16#34d2# => X"a9720000",
		16#34d3# => X"a4500001",
		16#34d4# => X"a86e0000",
		16#34d5# => X"a88d0000",
		16#34d6# => X"bc020000",
		16#34d7# => X"10000006",
		16#34d8# => X"ba100081",
		16#34d9# => X"84b40000",
		16#34da# => X"84d40004",
		16#34db# => X"07ffe4fe",
		16#34dc# => X"9f5a0001",
		16#34dd# => X"a9cb0000",
		16#34de# => X"a9ac0000",
		16#34df# => X"bc300000",
		16#34e0# => X"13fffff3",
		16#34e1# => X"9e940008",
		16#34e2# => X"aa4b0000",
		16#34e3# => X"03fffd4e",
		16#34e4# => X"d401602c",
		16#34e5# => X"18c00001",
		16#34e6# => X"9c84ffff",
		16#34e7# => X"a8c64118",
		16#34e8# => X"b9840003",
		16#34e9# => X"aaee0000",
		16#34ea# => X"aada0000",
		16#34eb# => X"e18c3000",
		16#34ec# => X"d4012050",
		16#34ed# => X"e0b60004",
		16#34ee# => X"e0d70004",
		16#34ef# => X"846c0000",
		16#34f0# => X"848c0004",
		16#34f1# => X"07ffe4e8",
		16#34f2# => X"aa920000",
		16#34f3# => X"8461002c",
		16#34f4# => X"84e10020",
		16#34f5# => X"aaa30000",
		16#34f6# => X"9ce70001",
		16#34f7# => X"e0740004",
		16#34f8# => X"e0950004",
		16#34f9# => X"d4013828",
		16#34fa# => X"d4016060",
		16#34fb# => X"07ffe849",
		16#34fc# => X"d4015854",
		16#34fd# => X"a86b0000",
		16#34fe# => X"07ffe7c1",
		16#34ff# => X"a9cb0000",
		16#3500# => X"85e1002c",
		16#3501# => X"e0ab0004",
		16#3502# => X"e0cc0004",
		16#3503# => X"aaaf0000",
		16#3504# => X"e0740004",
		16#3505# => X"e0950004",
		16#3506# => X"07ffe4b1",
		16#3507# => X"15000000",
		16#3508# => X"9dae0030",
		16#3509# => X"84610020",
		16#350a# => X"8441004c",
		16#350b# => X"d8036800",
		16#350c# => X"aacb0000",
		16#350d# => X"bc220001",
		16#350e# => X"0c00002a",
		16#350f# => X"aa8c0000",
		16#3510# => X"84c10020",
		16#3511# => X"84e1004c",
		16#3512# => X"87410028",
		16#3513# => X"e2463800",
		16#3514# => X"a9760000",
		16#3515# => X"18400001",
		16#3516# => X"a86b0000",
		16#3517# => X"a84240b0",
		16#3518# => X"84a20000",
		16#3519# => X"84c20004",
		16#351a# => X"07ffe4bf",
		16#351b# => X"a88c0000",
		16#351c# => X"aa0b0000",
		16#351d# => X"a88c0000",
		16#351e# => X"a8700000",
		16#351f# => X"07ffe825",
		16#3520# => X"a9cc0000",
		16#3521# => X"a86b0000",
		16#3522# => X"07ffe79d",
		16#3523# => X"aa8b0000",
		16#3524# => X"a8500000",
		16#3525# => X"a86e0000",
		16#3526# => X"e0ab0004",
		16#3527# => X"e0cc0004",
		16#3528# => X"e0830004",
		16#3529# => X"e0620004",
		16#352a# => X"07ffe48d",
		16#352b# => X"15000000",
		16#352c# => X"9c740030",
		16#352d# => X"d81a1800",
		16#352e# => X"9f5a0001",
		16#352f# => X"e43a9000",
		16#3530# => X"13ffffe6",
		16#3531# => X"18400001",
		16#3532# => X"84610028",
		16#3533# => X"84810050",
		16#3534# => X"aacb0000",
		16#3535# => X"e0632000",
		16#3536# => X"aa8c0000",
		16#3537# => X"d4011828",
		16#3538# => X"85a10054",
		16#3539# => X"84610060",
		16#353a# => X"19c00001",
		16#353b# => X"a9ed0000",
		16#353c# => X"aa030000",
		16#353d# => X"a9ce40c8",
		16#353e# => X"e06f0004",
		16#353f# => X"e0900004",
		16#3540# => X"84ae0000",
		16#3541# => X"84ce0004",
		16#3542# => X"07ffe456",
		16#3543# => X"aa140000",
		16#3544# => X"a9f60000",
		16#3545# => X"e0ab0004",
		16#3546# => X"e0cc0004",
		16#3547# => X"e06f0004",
		16#3548# => X"e0900004",
		16#3549# => X"07ffe6e2",
		16#354a# => X"15000000",
		16#354b# => X"bd4b0000",
		16#354c# => X"13fffc60",
		16#354d# => X"84610028",
		16#354e# => X"85810060",
		16#354f# => X"84410054",
		16#3550# => X"aa0c0000",
		16#3551# => X"a9e20000",
		16#3552# => X"846e0000",
		16#3553# => X"848e0004",
		16#3554# => X"e0af0004",
		16#3555# => X"e0d00004",
		16#3556# => X"07ffe461",
		16#3557# => X"a9d60000",
		16#3558# => X"a9f40000",
		16#3559# => X"e0ab0004",
		16#355a# => X"e0cc0004",
		16#355b# => X"e06e0004",
		16#355c# => X"e08f0004",
		16#355d# => X"07ffe70a",
		16#355e# => X"15000000",
		16#355f# => X"bd8b0000",
		16#3560# => X"0ffffb81",
		16#3561# => X"84c10008",
		16#3562# => X"00000003",
		16#3563# => X"84810028",
		16#3564# => X"a8820000",
		16#3565# => X"9c44ffff",
		16#3566# => X"90620000",
		16#3567# => X"bc030030",
		16#3568# => X"13fffffc",
		16#3569# => X"15000000",
		16#356a# => X"d4012028",
		16#356b# => X"8481005c",
		16#356c# => X"03fffd5a",
		16#356d# => X"d4012008",
		16#356e# => X"9c800000",
		16#356f# => X"03fffb4f",
		16#3570# => X"d4012044",
		16#3571# => X"9cc00001",
		16#3572# => X"d4013044",
		16#3573# => X"84410018",
		16#3574# => X"bda20000",
		16#3575# => X"1000002c",
		16#3576# => X"aa220000",
		16#3577# => X"d4011038",
		16#3578# => X"03fffb4e",
		16#3579# => X"d401101c",
		16#357a# => X"9ce00000",
		16#357b# => X"03fffff8",
		16#357c# => X"d4013844",
		16#357d# => X"84610030",
		16#357e# => X"04000aad",
		16#357f# => X"a8820000",
		16#3580# => X"bd6b0000",
		16#3581# => X"13fffdd4",
		16#3582# => X"84c1001c",
		16#3583# => X"84e10008",
		16#3584# => X"a87e0000",
		16#3585# => X"84810030",
		16#3586# => X"9ce7ffff",
		16#3587# => X"9ca0000a",
		16#3588# => X"9cc00000",
		16#3589# => X"04000859",
		16#358a# => X"d4013808",
		16#358b# => X"84610038",
		16#358c# => X"84810044",
		16#358d# => X"d4015830",
		16#358e# => X"bc040000",
		16#358f# => X"13fffdc5",
		16#3590# => X"d401181c",
		16#3591# => X"a8920000",
		16#3592# => X"a87e0000",
		16#3593# => X"9ca0000a",
		16#3594# => X"0400084e",
		16#3595# => X"9cc00000",
		16#3596# => X"03fffdbe",
		16#3597# => X"aa4b0000",
		16#3598# => X"85820010",
		16#3599# => X"9d8c0004",
		16#359a# => X"b98c0002",
		16#359b# => X"e1826000",
		16#359c# => X"040008d6",
		16#359d# => X"846c0000",
		16#359e# => X"9da00020",
		16#359f# => X"03fffd92",
		16#35a0# => X"e1ad5802",
		16#35a1# => X"9c600001",
		16#35a2# => X"d4011838",
		16#35a3# => X"d401181c",
		16#35a4# => X"03fffc50",
		16#35a5# => X"d4011818",
		16#35a6# => X"bcb1000e",
		16#35a7# => X"10000003",
		16#35a8# => X"9d800001",
		16#35a9# => X"9d800000",
		16#35aa# => X"e1ce6003",
		16#35ab# => X"03fffc49",
		16#35ac# => X"d401881c",
		16#35ad# => X"84e10010",
		16#35ae# => X"e4278000",
		16#35af# => X"13fffd7f",
		16#35b0# => X"84610048",
		16#35b1# => X"1860000f",
		16#35b2# => X"a863ffff",
		16#35b3# => X"e19c1803",
		16#35b4# => X"bc2c0000",
		16#35b5# => X"13fffd78",
		16#35b6# => X"aa070000",
		16#35b7# => X"18807ff0",
		16#35b8# => X"e39c2003",
		16#35b9# => X"bc1c0000",
		16#35ba# => X"13fffd74",
		16#35bb# => X"84610048",
		16#35bc# => X"84c10034",
		16#35bd# => X"84e10024",
		16#35be# => X"9cc60001",
		16#35bf# => X"9ce70001",
		16#35c0# => X"d4013034",
		16#35c1# => X"d4013824",
		16#35c2# => X"03fffd6b",
		16#35c3# => X"9e000001",
		16#35c4# => X"10000006",
		16#35c5# => X"a8920000",
		16#35c6# => X"a87e0000",
		16#35c7# => X"04000a05",
		16#35c8# => X"a8ae0000",
		16#35c9# => X"aa4b0000",
		16#35ca# => X"bc100000",
		16#35cb# => X"0c0000bd",
		16#35cc# => X"aa920000",
		16#35cd# => X"9f400001",
		16#35ce# => X"84c10010",
		16#35cf# => X"84810020",
		16#35d0# => X"e386d003",
		16#35d1# => X"d4012028",
		16#35d2# => X"d401e018",
		16#35d3# => X"a9d20000",
		16#35d4# => X"ab9a0000",
		16#35d5# => X"87010030",
		16#35d6# => X"ab440000",
		16#35d7# => X"a8780000",
		16#35d8# => X"a8820000",
		16#35d9# => X"07fff945",
		16#35da# => X"9ec00001",
		16#35db# => X"a8780000",
		16#35dc# => X"a88e0000",
		16#35dd# => X"9d6b0030",
		16#35de# => X"04000a4d",
		16#35df# => X"d4015810",
		16#35e0# => X"a87e0000",
		16#35e1# => X"a8820000",
		16#35e2# => X"a8b40000",
		16#35e3# => X"04000a63",
		16#35e4# => X"aa0b0000",
		16#35e5# => X"846b000c",
		16#35e6# => X"bc230000",
		16#35e7# => X"0c000035",
		16#35e8# => X"aa4b0000",
		16#35e9# => X"a87e0000",
		16#35ea# => X"040007ec",
		16#35eb# => X"a8920000",
		16#35ec# => X"84e10000",
		16#35ed# => X"e0763804",
		16#35ee# => X"bc230000",
		16#35ef# => X"10000006",
		16#35f0# => X"bd900000",
		16#35f1# => X"84610018",
		16#35f2# => X"bc230000",
		16#35f3# => X"0c0000c4",
		16#35f4# => X"bd900000",
		16#35f5# => X"10000067",
		16#35f6# => X"84c10000",
		16#35f7# => X"e2103004",
		16#35f8# => X"bc300000",
		16#35f9# => X"10000006",
		16#35fa# => X"bdb60000",
		16#35fb# => X"84e10018",
		16#35fc# => X"bc270000",
		16#35fd# => X"0c00005f",
		16#35fe# => X"bdb60000",
		16#35ff# => X"0c0000a3",
		16#3600# => X"84610010",
		16#3601# => X"d81a1800",
		16#3602# => X"8481001c",
		16#3603# => X"e41c2000",
		16#3604# => X"10000099",
		16#3605# => X"9f5a0001",
		16#3606# => X"a8980000",
		16#3607# => X"a87e0000",
		16#3608# => X"9ca0000a",
		16#3609# => X"040007d9",
		16#360a# => X"9cc00000",
		16#360b# => X"e42ea000",
		16#360c# => X"0c000015",
		16#360d# => X"ab0b0000",
		16#360e# => X"a88e0000",
		16#360f# => X"9ca0000a",
		16#3610# => X"9cc00000",
		16#3611# => X"a87e0000",
		16#3612# => X"040007d0",
		16#3613# => X"9f9c0001",
		16#3614# => X"a8940000",
		16#3615# => X"a87e0000",
		16#3616# => X"9ca0000a",
		16#3617# => X"9cc00000",
		16#3618# => X"040007ca",
		16#3619# => X"a9cb0000",
		16#361a# => X"03ffffbd",
		16#361b# => X"aa8b0000",
		16#361c# => X"a8780000",
		16#361d# => X"04000a0e",
		16#361e# => X"a88b0000",
		16#361f# => X"03ffffca",
		16#3620# => X"aacb0000",
		16#3621# => X"a88e0000",
		16#3622# => X"a87e0000",
		16#3623# => X"9ca0000a",
		16#3624# => X"9cc00000",
		16#3625# => X"040007bd",
		16#3626# => X"9f9c0001",
		16#3627# => X"a9cb0000",
		16#3628# => X"03ffffaf",
		16#3629# => X"aa8b0000",
		16#362a# => X"03fffc9c",
		16#362b# => X"d401b028",
		16#362c# => X"a87e0000",
		16#362d# => X"84810030",
		16#362e# => X"04000946",
		16#362f# => X"84a10040",
		16#3630# => X"03fffced",
		16#3631# => X"d4015830",
		16#3632# => X"84610048",
		16#3633# => X"e1901002",
		16#3634# => X"9e000000",
		16#3635# => X"e0636000",
		16#3636# => X"e0426000",
		16#3637# => X"d4011848",
		16#3638# => X"03fffcaa",
		16#3639# => X"d4011040",
		16#363a# => X"84810030",
		16#363b# => X"04000939",
		16#363c# => X"a8b00000",
		16#363d# => X"03fffce0",
		16#363e# => X"d4015830",
		16#363f# => X"9c400000",
		16#3640# => X"03fffc72",
		16#3641# => X"aa420000",
		16#3642# => X"84810058",
		16#3643# => X"bc040000",
		16#3644# => X"10000054",
		16#3645# => X"9c400036",
		16#3646# => X"9dad0433",
		16#3647# => X"86010040",
		16#3648# => X"03fffca0",
		16#3649# => X"85c10034",
		16#364a# => X"9cc60001",
		16#364b# => X"d4011828",
		16#364c# => X"b8c60018",
		16#364d# => X"8461005c",
		16#364e# => X"d4012020",
		16#364f# => X"b8c60098",
		16#3650# => X"d4011808",
		16#3651# => X"03fffc75",
		16#3652# => X"d8023000",
		16#3653# => X"84810020",
		16#3654# => X"03fffb5b",
		16#3655# => X"87c10060",
		16#3656# => X"87c10060",
		16#3657# => X"03fffa89",
		16#3658# => X"87810064",
		16#3659# => X"9da00000",
		16#365a# => X"03fffc8e",
		16#365b# => X"e1c62002",
		16#365c# => X"d401c030",
		16#365d# => X"d401d028",
		16#365e# => X"bdb60000",
		16#365f# => X"1000000f",
		16#3660# => X"86010010",
		16#3661# => X"9ca00001",
		16#3662# => X"a87e0000",
		16#3663# => X"04000969",
		16#3664# => X"a8980000",
		16#3665# => X"a8820000",
		16#3666# => X"a86b0000",
		16#3667# => X"040009c4",
		16#3668# => X"d4015830",
		16#3669# => X"bd4b0000",
		16#366a# => X"0c00005d",
		16#366b# => X"bc100039",
		16#366c# => X"10000042",
		16#366d# => X"9e100001",
		16#366e# => X"84610028",
		16#366f# => X"aa540000",
		16#3670# => X"d8038000",
		16#3671# => X"9c630001",
		16#3672# => X"03fffc46",
		16#3673# => X"d4011828",
		16#3674# => X"10000009",
		16#3675# => X"84a10028",
		16#3676# => X"a6100001",
		16#3677# => X"bc300000",
		16#3678# => X"13fffe19",
		16#3679# => X"84610028",
		16#367a# => X"00000004",
		16#367b# => X"9c65ffff",
		16#367c# => X"a8a30000",
		16#367d# => X"9c65ffff",
		16#367e# => X"90830000",
		16#367f# => X"bc040030",
		16#3680# => X"13fffffc",
		16#3681# => X"15000000",
		16#3682# => X"03fffc36",
		16#3683# => X"d4012828",
		16#3684# => X"9ce70001",
		16#3685# => X"d4011828",
		16#3686# => X"03fffc32",
		16#3687# => X"d8063800",
		16#3688# => X"a87e0000",
		16#3689# => X"04000720",
		16#368a# => X"84920004",
		16#368b# => X"84f20010",
		16#368c# => X"9c6b000c",
		16#368d# => X"9ce70002",
		16#368e# => X"9c92000c",
		16#368f# => X"b8a70002",
		16#3690# => X"04000626",
		16#3691# => X"a9cb0000",
		16#3692# => X"a87e0000",
		16#3693# => X"a88e0000",
		16#3694# => X"04000938",
		16#3695# => X"9ca00001",
		16#3696# => X"03ffff37",
		16#3697# => X"aa8b0000",
		16#3698# => X"85a1006c",
		16#3699# => X"86010040",
		16#369a# => X"e1a26802",
		16#369b# => X"03fffc4d",
		16#369c# => X"85c10034",
		16#369d# => X"86010010",
		16#369e# => X"d401c030",
		16#369f# => X"d401d028",
		16#36a0# => X"03fffde5",
		16#36a1# => X"aa540000",
		16#36a2# => X"86010010",
		16#36a3# => X"d401c030",
		16#36a4# => X"bc300039",
		16#36a5# => X"0c000009",
		16#36a6# => X"d401d028",
		16#36a7# => X"84e10028",
		16#36a8# => X"9e100001",
		16#36a9# => X"aa540000",
		16#36aa# => X"d8078000",
		16#36ab# => X"9ce70001",
		16#36ac# => X"03fffc0c",
		16#36ad# => X"d4013828",
		16#36ae# => X"84810028",
		16#36af# => X"9cc00039",
		16#36b0# => X"aa540000",
		16#36b1# => X"d8043000",
		16#36b2# => X"9c840001",
		16#36b3# => X"d4012028",
		16#36b4# => X"a8640000",
		16#36b5# => X"03fffddf",
		16#36b6# => X"84810020",
		16#36b7# => X"d401c030",
		16#36b8# => X"d401d028",
		16#36b9# => X"ab100000",
		16#36ba# => X"86010010",
		16#36bb# => X"bc100039",
		16#36bc# => X"13fffff2",
		16#36bd# => X"bdb80000",
		16#36be# => X"10000003",
		16#36bf# => X"15000000",
		16#36c0# => X"9e100001",
		16#36c1# => X"84810028",
		16#36c2# => X"aa540000",
		16#36c3# => X"d8048000",
		16#36c4# => X"9c840001",
		16#36c5# => X"03fffbf3",
		16#36c6# => X"d4012028",
		16#36c7# => X"bc2b0000",
		16#36c8# => X"13ffffa7",
		16#36c9# => X"84610028",
		16#36ca# => X"a4700001",
		16#36cb# => X"bc030000",
		16#36cc# => X"13ffffa3",
		16#36cd# => X"84610028",
		16#36ce# => X"03ffff9e",
		16#36cf# => X"bc100039",
		16#36d0# => X"8481005c",
		16#36d1# => X"03fffbf5",
		16#36d2# => X"d4012008",
		16#36d3# => X"8461001c",
		16#36d4# => X"bca3000e",
		16#36d5# => X"10000003",
		16#36d6# => X"9c400001",
		16#36d7# => X"9c400000",
		16#36d8# => X"e1ce1003",
		16#36d9# => X"03fffb1d",
		16#36da# => X"9c400000",
		16#36db# => X"bc0c0004",
		16#36dc# => X"13fffc63",
		16#36dd# => X"84810034",
		16#36de# => X"03fffc59",
		16#36df# => X"9d8c001c",
		16#36e0# => X"d7e117ec",
		16#36e1# => X"d7e197f8",
		16#36e2# => X"d7e14ffc",
		16#36e3# => X"d7e177f0",
		16#36e4# => X"d7e187f4",
		16#36e5# => X"aa430000",
		16#36e6# => X"9c21ffec",
		16#36e7# => X"bc030000",
		16#36e8# => X"10000006",
		16#36e9# => X"a8440000",
		16#36ea# => X"84830038",
		16#36eb# => X"bc240000",
		16#36ec# => X"0c00007b",
		16#36ed# => X"15000000",
		16#36ee# => X"9962000c",
		16#36ef# => X"bc0b0000",
		16#36f0# => X"10000048",
		16#36f1# => X"a88b0000",
		16#36f2# => X"a46b0008",
		16#36f3# => X"bc230000",
		16#36f4# => X"1000004b",
		16#36f5# => X"15000000",
		16#36f6# => X"a88b0800",
		16#36f7# => X"84a20004",
		16#36f8# => X"bd450000",
		16#36f9# => X"0c000086",
		16#36fa# => X"dc02200c",
		16#36fb# => X"84e20028",
		16#36fc# => X"bc070000",
		16#36fd# => X"1000003b",
		16#36fe# => X"a9670000",
		16#36ff# => X"a464ffff",
		16#3700# => X"9c800000",
		16#3701# => X"85d20000",
		16#3702# => X"a4a31000",
		16#3703# => X"e4052000",
		16#3704# => X"10000069",
		16#3705# => X"d4122000",
		16#3706# => X"84a20050",
		16#3707# => X"a4630004",
		16#3708# => X"bc030000",
		16#3709# => X"1000000a",
		16#370a# => X"a8720000",
		16#370b# => X"84820004",
		16#370c# => X"84620030",
		16#370d# => X"bc030000",
		16#370e# => X"10000004",
		16#370f# => X"e0a52002",
		16#3710# => X"8462003c",
		16#3711# => X"e0a51802",
		16#3712# => X"a8720000",
		16#3713# => X"8482001c",
		16#3714# => X"48003800",
		16#3715# => X"9cc00000",
		16#3716# => X"bc2bffff",
		16#3717# => X"0c00006e",
		16#3718# => X"15000000",
		16#3719# => X"9462000c",
		16#371a# => X"9ca0f7ff",
		16#371b# => X"84820010",
		16#371c# => X"e0632803",
		16#371d# => X"9ca00000",
		16#371e# => X"b8630010",
		16#371f# => X"d4022000",
		16#3720# => X"d4022804",
		16#3721# => X"b8630090",
		16#3722# => X"a4831000",
		16#3723# => X"e4042800",
		16#3724# => X"10000006",
		16#3725# => X"dc02180c",
		16#3726# => X"bc2bffff",
		16#3727# => X"0c00006a",
		16#3728# => X"15000000",
		16#3729# => X"d4025850",
		16#372a# => X"84820030",
		16#372b# => X"d4127000",
		16#372c# => X"bc040000",
		16#372d# => X"1000000b",
		16#372e# => X"a9640000",
		16#372f# => X"9c620040",
		16#3730# => X"e4041800",
		16#3731# => X"10000005",
		16#3732# => X"9c600000",
		16#3733# => X"040001dc",
		16#3734# => X"a8720000",
		16#3735# => X"9c600000",
		16#3736# => X"d4021830",
		16#3737# => X"a9630000",
		16#3738# => X"9c210014",
		16#3739# => X"8521fffc",
		16#373a# => X"8441ffec",
		16#373b# => X"85c1fff0",
		16#373c# => X"8601fff4",
		16#373d# => X"44004800",
		16#373e# => X"8641fff8",
		16#373f# => X"85c20010",
		16#3740# => X"bc0e0000",
		16#3741# => X"13fffff7",
		16#3742# => X"a96e0000",
		16#3743# => X"86020000",
		16#3744# => X"a4840003",
		16#3745# => X"9c600000",
		16#3746# => X"d4027000",
		16#3747# => X"e4241800",
		16#3748# => X"0c000023",
		16#3749# => X"e2107002",
		16#374a# => X"9d600000",
		16#374b# => X"e5b05800",
		16#374c# => X"0c000007",
		16#374d# => X"d4021808",
		16#374e# => X"03ffffeb",
		16#374f# => X"9c210014",
		16#3750# => X"bdb00000",
		16#3751# => X"10000026",
		16#3752# => X"e1ce5800",
		16#3753# => X"a8d00000",
		16#3754# => X"a8ae0000",
		16#3755# => X"85620024",
		16#3756# => X"a8720000",
		16#3757# => X"48005800",
		16#3758# => X"8482001c",
		16#3759# => X"bd4b0000",
		16#375a# => X"13fffff6",
		16#375b# => X"e2105802",
		16#375c# => X"9462000c",
		16#375d# => X"a8630040",
		16#375e# => X"9d60ffff",
		16#375f# => X"dc02180c",
		16#3760# => X"9c210014",
		16#3761# => X"8521fffc",
		16#3762# => X"8441ffec",
		16#3763# => X"85c1fff0",
		16#3764# => X"8601fff4",
		16#3765# => X"44004800",
		16#3766# => X"8641fff8",
		16#3767# => X"04000087",
		16#3768# => X"15000000",
		16#3769# => X"03ffff86",
		16#376a# => X"9962000c",
		16#376b# => X"03ffffdf",
		16#376c# => X"84620014",
		16#376d# => X"a8720000",
		16#376e# => X"8482001c",
		16#376f# => X"48003800",
		16#3770# => X"9cc00001",
		16#3771# => X"bc2bffff",
		16#3772# => X"0c000025",
		16#3773# => X"a8ab0000",
		16#3774# => X"9462000c",
		16#3775# => X"03ffff92",
		16#3776# => X"84e20028",
		16#3777# => X"9c210014",
		16#3778# => X"9d600000",
		16#3779# => X"8521fffc",
		16#377a# => X"8441ffec",
		16#377b# => X"85c1fff0",
		16#377c# => X"8601fff4",
		16#377d# => X"44004800",
		16#377e# => X"8641fff8",
		16#377f# => X"84a2003c",
		16#3780# => X"bda50000",
		16#3781# => X"0fffff7a",
		16#3782# => X"a9630000",
		16#3783# => X"03ffffb6",
		16#3784# => X"9c210014",
		16#3785# => X"84720000",
		16#3786# => X"bc030000",
		16#3787# => X"13ffff92",
		16#3788# => X"bc03001d",
		16#3789# => X"13ffff90",
		16#378a# => X"bc230016",
		16#378b# => X"0fffff8e",
		16#378c# => X"15000000",
		16#378d# => X"9462000c",
		16#378e# => X"a8630040",
		16#378f# => X"03ffffa9",
		16#3790# => X"dc02180c",
		16#3791# => X"84720000",
		16#3792# => X"e4232800",
		16#3793# => X"13ffff97",
		16#3794# => X"15000000",
		16#3795# => X"03ffff95",
		16#3796# => X"d4025850",
		16#3797# => X"84720000",
		16#3798# => X"bc230000",
		16#3799# => X"0fffffdb",
		16#379a# => X"ac830016",
		16#379b# => X"e0c02002",
		16#379c# => X"e0862004",
		16#379d# => X"bd640000",
		16#379e# => X"10000007",
		16#379f# => X"ac63001d",
		16#37a0# => X"e0801802",
		16#37a1# => X"e0641804",
		16#37a2# => X"bd830000",
		16#37a3# => X"10000005",
		16#37a4# => X"15000000",
		16#37a5# => X"d4127000",
		16#37a6# => X"03ffff92",
		16#37a7# => X"9d600000",
		16#37a8# => X"9462000c",
		16#37a9# => X"a8630040",
		16#37aa# => X"03ffff8e",
		16#37ab# => X"dc02180c",
		16#37ac# => X"d7e14ffc",
		16#37ad# => X"bc230000",
		16#37ae# => X"0c00000a",
		16#37af# => X"9c21fffc",
		16#37b0# => X"a8830000",
		16#37b1# => X"18600001",
		16#37b2# => X"a86363e0",
		16#37b3# => X"84630000",
		16#37b4# => X"9c210004",
		16#37b5# => X"8521fffc",
		16#37b6# => X"03ffff2a",
		16#37b7# => X"15000000",
		16#37b8# => X"18600001",
		16#37b9# => X"18800000",
		16#37ba# => X"a8633ea0",
		16#37bb# => X"9c210004",
		16#37bc# => X"a884db80",
		16#37bd# => X"8521fffc",
		16#37be# => X"000003c0",
		16#37bf# => X"84630000",
		16#37c0# => X"44004800",
		16#37c1# => X"9d600000",
		16#37c2# => X"44004800",
		16#37c3# => X"9d600000",
		16#37c4# => X"d7e14ffc",
		16#37c5# => X"9c21fffc",
		16#37c6# => X"18800001",
		16#37c7# => X"9c210004",
		16#37c8# => X"8521fffc",
		16#37c9# => X"00000383",
		16#37ca# => X"a88429e4",
		16#37cb# => X"d7e177f4",
		16#37cc# => X"9dc00068",
		16#37cd# => X"d7e117f0",
		16#37ce# => X"e1c47306",
		16#37cf# => X"d7e187f8",
		16#37d0# => X"d7e14ffc",
		16#37d1# => X"aa040000",
		16#37d2# => X"9c21fff0",
		16#37d3# => X"07ffe687",
		16#37d4# => X"9c8e000c",
		16#37d5# => X"bc0b0000",
		16#37d6# => X"10000009",
		16#37d7# => X"a84b0000",
		16#37d8# => X"9c6b000c",
		16#37d9# => X"9c800000",
		16#37da# => X"d40b8004",
		16#37db# => X"d40b2000",
		16#37dc# => X"d40b1808",
		16#37dd# => X"0400057c",
		16#37de# => X"a8ae0000",
		16#37df# => X"9c210010",
		16#37e0# => X"a9620000",
		16#37e1# => X"8521fffc",
		16#37e2# => X"8441fff0",
		16#37e3# => X"85c1fff4",
		16#37e4# => X"44004800",
		16#37e5# => X"8601fff8",
		16#37e6# => X"d7e14ffc",
		16#37e7# => X"18600001",
		16#37e8# => X"9c21fffc",
		16#37e9# => X"a8633ea0",
		16#37ea# => X"9c210004",
		16#37eb# => X"8521fffc",
		16#37ec# => X"03ffffd8",
		16#37ed# => X"84630000",
		16#37ee# => X"d7e117d8",
		16#37ef# => X"d7e197e4",
		16#37f0# => X"d7e14ffc",
		16#37f1# => X"d7e177dc",
		16#37f2# => X"d7e187e0",
		16#37f3# => X"d7e1a7e8",
		16#37f4# => X"d7e1b7ec",
		16#37f5# => X"d7e1c7f0",
		16#37f6# => X"d7e1d7f4",
		16#37f7# => X"d7e1e7f8",
		16#37f8# => X"84430038",
		16#37f9# => X"9c21ffd8",
		16#37fa# => X"bc220000",
		16#37fb# => X"10000051",
		16#37fc# => X"aa430000",
		16#37fd# => X"18800000",
		16#37fe# => X"9f800001",
		16#37ff# => X"a884df10",
		16#3800# => X"9c6302ec",
		16#3801# => X"d412203c",
		16#3802# => X"9c800003",
		16#3803# => X"85d20004",
		16#3804# => X"9cc00004",
		16#3805# => X"d41222e4",
		16#3806# => X"d4121ae8",
		16#3807# => X"d412e038",
		16#3808# => X"d41212e0",
		16#3809# => X"9c6e005c",
		16#380a# => X"dc0e300c",
		16#380b# => X"a8820000",
		16#380c# => X"9ca00008",
		16#380d# => X"d40e1000",
		16#380e# => X"d40e1004",
		16#380f# => X"d40e1008",
		16#3810# => X"d40e1064",
		16#3811# => X"dc0e100e",
		16#3812# => X"d40e1010",
		16#3813# => X"d40e1014",
		16#3814# => X"d40e1018",
		16#3815# => X"1b400001",
		16#3816# => X"1b000001",
		16#3817# => X"1ac00001",
		16#3818# => X"04000541",
		16#3819# => X"1a800001",
		16#381a# => X"ab5a135c",
		16#381b# => X"86120008",
		16#381c# => X"ab1813c0",
		16#381d# => X"aad61444",
		16#381e# => X"aa9414a4",
		16#381f# => X"9cc00009",
		16#3820# => X"9c70005c",
		16#3821# => X"a8820000",
		16#3822# => X"9ca00008",
		16#3823# => X"d40e701c",
		16#3824# => X"d40ed020",
		16#3825# => X"d40ec024",
		16#3826# => X"d40eb028",
		16#3827# => X"d40ea02c",
		16#3828# => X"dc10300c",
		16#3829# => X"d4101000",
		16#382a# => X"d4101004",
		16#382b# => X"d4101008",
		16#382c# => X"d4101064",
		16#382d# => X"dc10e00e",
		16#382e# => X"d4101010",
		16#382f# => X"d4101014",
		16#3830# => X"04000529",
		16#3831# => X"d4101018",
		16#3832# => X"9c600012",
		16#3833# => X"85d2000c",
		16#3834# => X"9cc00002",
		16#3835# => X"dc0e180c",
		16#3836# => X"d410801c",
		16#3837# => X"d410d020",
		16#3838# => X"d410c024",
		16#3839# => X"d410b028",
		16#383a# => X"d410a02c",
		16#383b# => X"d40e1000",
		16#383c# => X"d40e1004",
		16#383d# => X"d40e1008",
		16#383e# => X"d40e1064",
		16#383f# => X"dc0e300e",
		16#3840# => X"d40e1010",
		16#3841# => X"d40e1014",
		16#3842# => X"d40e1018",
		16#3843# => X"9c6e005c",
		16#3844# => X"a8820000",
		16#3845# => X"04000514",
		16#3846# => X"9ca00008",
		16#3847# => X"d40e701c",
		16#3848# => X"d40ed020",
		16#3849# => X"d40ec024",
		16#384a# => X"d40eb028",
		16#384b# => X"d40ea02c",
		16#384c# => X"9c210028",
		16#384d# => X"8521fffc",
		16#384e# => X"8441ffd8",
		16#384f# => X"85c1ffdc",
		16#3850# => X"8601ffe0",
		16#3851# => X"8641ffe4",
		16#3852# => X"8681ffe8",
		16#3853# => X"86c1ffec",
		16#3854# => X"8701fff0",
		16#3855# => X"8741fff4",
		16#3856# => X"44004800",
		16#3857# => X"8781fff8",
		16#3858# => X"d7e117f0",
		16#3859# => X"18400001",
		16#385a# => X"d7e177f4",
		16#385b# => X"a8423ea0",
		16#385c# => X"d7e187f8",
		16#385d# => X"85c20000",
		16#385e# => X"d7e14ffc",
		16#385f# => X"844e0038",
		16#3860# => X"9c21fff0",
		16#3861# => X"bc220000",
		16#3862# => X"0c000033",
		16#3863# => X"aa030000",
		16#3864# => X"9dce02e0",
		16#3865# => X"848e0004",
		16#3866# => X"9c84ffff",
		16#3867# => X"bd840000",
		16#3868# => X"0c000007",
		16#3869# => X"844e0008",
		16#386a# => X"00000026",
		16#386b# => X"856e0000",
		16#386c# => X"bd640000",
		16#386d# => X"0c000022",
		16#386e# => X"9c420068",
		16#386f# => X"98a2000c",
		16#3870# => X"bc050000",
		16#3871# => X"0ffffffb",
		16#3872# => X"9c84ffff",
		16#3873# => X"9c60ffff",
		16#3874# => X"9c800000",
		16#3875# => X"dc02180e",
		16#3876# => X"9c600001",
		16#3877# => X"9ca00008",
		16#3878# => X"dc02180c",
		16#3879# => X"9c600000",
		16#387a# => X"d4021864",
		16#387b# => X"d4021800",
		16#387c# => X"d4021808",
		16#387d# => X"d4021804",
		16#387e# => X"d4021810",
		16#387f# => X"d4021814",
		16#3880# => X"d4021818",
		16#3881# => X"040004d8",
		16#3882# => X"9c62005c",
		16#3883# => X"9c600000",
		16#3884# => X"d4021830",
		16#3885# => X"d4021834",
		16#3886# => X"d4021844",
		16#3887# => X"d4021848",
		16#3888# => X"9c210010",
		16#3889# => X"a9620000",
		16#388a# => X"8521fffc",
		16#388b# => X"8441fff0",
		16#388c# => X"85c1fff4",
		16#388d# => X"44004800",
		16#388e# => X"8601fff8",
		16#388f# => X"856e0000",
		16#3890# => X"bc2b0000",
		16#3891# => X"0c000008",
		16#3892# => X"15000000",
		16#3893# => X"03ffffd2",
		16#3894# => X"a9cb0000",
		16#3895# => X"07ffff59",
		16#3896# => X"a86e0000",
		16#3897# => X"03ffffce",
		16#3898# => X"9dce02e0",
		16#3899# => X"a8700000",
		16#389a# => X"07ffff31",
		16#389b# => X"9c800004",
		16#389c# => X"bc0b0000",
		16#389d# => X"0ffffff6",
		16#389e# => X"d40e5800",
		16#389f# => X"9c60000c",
		16#38a0# => X"a84b0000",
		16#38a1# => X"03ffffe7",
		16#38a2# => X"d4101800",
		16#38a3# => X"44004800",
		16#38a4# => X"15000000",
		16#38a5# => X"44004800",
		16#38a6# => X"15000000",
		16#38a7# => X"44004800",
		16#38a8# => X"15000000",
		16#38a9# => X"44004800",
		16#38aa# => X"15000000",
		16#38ab# => X"18600001",
		16#38ac# => X"d7e14ffc",
		16#38ad# => X"a86363e0",
		16#38ae# => X"9c21fffc",
		16#38af# => X"18800000",
		16#38b0# => X"84630000",
		16#38b1# => X"9c210004",
		16#38b2# => X"8521fffc",
		16#38b3# => X"00000299",
		16#38b4# => X"a884df00",
		16#38b5# => X"18600001",
		16#38b6# => X"d7e14ffc",
		16#38b7# => X"a86363e0",
		16#38b8# => X"9c21fffc",
		16#38b9# => X"18800000",
		16#38ba# => X"84630000",
		16#38bb# => X"9c210004",
		16#38bc# => X"8521fffc",
		16#38bd# => X"0000028f",
		16#38be# => X"a884df08",
		16#38bf# => X"d7e117ec",
		16#38c0# => X"18400001",
		16#38c1# => X"d7e177f0",
		16#38c2# => X"d7e187f4",
		16#38c3# => X"d7e197f8",
		16#38c4# => X"d7e14ffc",
		16#38c5# => X"9c21ffec",
		16#38c6# => X"a8426808",
		16#38c7# => X"aa440000",
		16#38c8# => X"07ffe7e2",
		16#38c9# => X"a9c30000",
		16#38ca# => X"84620008",
		16#38cb# => X"86030004",
		16#38cc# => X"9c60fffc",
		16#38cd# => X"e2101803",
		16#38ce# => X"9c700fef",
		16#38cf# => X"e2439002",
		16#38d0# => X"9c60f000",
		16#38d1# => X"e2521803",
		16#38d2# => X"e2521800",
		16#38d3# => X"bd520fff",
		16#38d4# => X"0c000009",
		16#38d5# => X"a86e0000",
		16#38d6# => X"07ffec6a",
		16#38d7# => X"9c800000",
		16#38d8# => X"84620008",
		16#38d9# => X"e0638000",
		16#38da# => X"e40b1800",
		16#38db# => X"1000000c",
		16#38dc# => X"a86e0000",
		16#38dd# => X"07ffe7cf",
		16#38de# => X"a86e0000",
		16#38df# => X"9c210014",
		16#38e0# => X"9d600000",
		16#38e1# => X"8521fffc",
		16#38e2# => X"8441ffec",
		16#38e3# => X"85c1fff0",
		16#38e4# => X"8601fff4",
		16#38e5# => X"44004800",
		16#38e6# => X"8641fff8",
		16#38e7# => X"07ffec59",
		16#38e8# => X"e0809002",
		16#38e9# => X"bc2bffff",
		16#38ea# => X"0c000014",
		16#38eb# => X"18800001",
		16#38ec# => X"e2109002",
		16#38ed# => X"a8847a84",
		16#38ee# => X"84420008",
		16#38ef# => X"84640000",
		16#38f0# => X"aa100001",
		16#38f1# => X"e2439002",
		16#38f2# => X"d4028004",
		16#38f3# => X"a86e0000",
		16#38f4# => X"07ffe7b8",
		16#38f5# => X"d4049000",
		16#38f6# => X"9c210014",
		16#38f7# => X"9d600001",
		16#38f8# => X"8521fffc",
		16#38f9# => X"8441ffec",
		16#38fa# => X"85c1fff0",
		16#38fb# => X"8601fff4",
		16#38fc# => X"44004800",
		16#38fd# => X"8641fff8",
		16#38fe# => X"a86e0000",
		16#38ff# => X"07ffec41",
		16#3900# => X"9c800000",
		16#3901# => X"84420008",
		16#3902# => X"e06b1002",
		16#3903# => X"bda3000f",
		16#3904# => X"13ffffd9",
		16#3905# => X"18800001",
		16#3906# => X"a8630001",
		16#3907# => X"a8846c14",
		16#3908# => X"d4021804",
		16#3909# => X"84840000",
		16#390a# => X"18400001",
		16#390b# => X"e16b2002",
		16#390c# => X"a8427a84",
		16#390d# => X"03ffffd0",
		16#390e# => X"d4025800",
		16#390f# => X"d7e117f4",
		16#3910# => X"d7e177f8",
		16#3911# => X"d7e14ffc",
		16#3912# => X"a9c40000",
		16#3913# => X"9c21fff4",
		16#3914# => X"bc040000",
		16#3915# => X"10000062",
		16#3916# => X"a8430000",
		16#3917# => X"07ffe793",
		16#3918# => X"15000000",
		16#3919# => X"9c8efff8",
		16#391a# => X"9c60fffe",
		16#391b# => X"18e00001",
		16#391c# => X"85040004",
		16#391d# => X"a8e76808",
		16#391e# => X"e0a81803",
		16#391f# => X"85670008",
		16#3920# => X"e0c42800",
		16#3921# => X"84660004",
		16#3922# => X"e42b3000",
		16#3923# => X"9d60fffc",
		16#3924# => X"0c00007c",
		16#3925# => X"e0635803",
		16#3926# => X"a5080001",
		16#3927# => X"9d600000",
		16#3928# => X"e4285800",
		16#3929# => X"1000000f",
		16#392a# => X"d4061804",
		16#392b# => X"85840000",
		16#392c# => X"19a00001",
		16#392d# => X"e0846002",
		16#392e# => X"e0a56000",
		16#392f# => X"a9ad6810",
		16#3930# => X"85840008",
		16#3931# => X"e40c6800",
		16#3932# => X"10000006",
		16#3933# => X"9d600001",
		16#3934# => X"85a4000c",
		16#3935# => X"a9680000",
		16#3936# => X"d40c680c",
		16#3937# => X"d40d6008",
		16#3938# => X"e1061800",
		16#3939# => X"85080004",
		16#393a# => X"a5080001",
		16#393b# => X"bc280000",
		16#393c# => X"10000008",
		16#393d# => X"bc2b0000",
		16#393e# => X"0c00003e",
		16#393f# => X"e0a51800",
		16#3940# => X"84660008",
		16#3941# => X"84c6000c",
		16#3942# => X"d403300c",
		16#3943# => X"d4061808",
		16#3944# => X"a8c50001",
		16#3945# => X"e0642800",
		16#3946# => X"d4043004",
		16#3947# => X"bc2b0000",
		16#3948# => X"10000029",
		16#3949# => X"d4032800",
		16#394a# => X"bc4501ff",
		16#394b# => X"0c000040",
		16#394c# => X"9cc00001",
		16#394d# => X"b8650049",
		16#394e# => X"bc430004",
		16#394f# => X"1000006b",
		16#3950# => X"bc430014",
		16#3951# => X"b9050046",
		16#3952# => X"9d080038",
		16#3953# => X"b8680003",
		16#3954# => X"19a00001",
		16#3955# => X"a9ad6808",
		16#3956# => X"e0636800",
		16#3957# => X"84c30008",
		16#3958# => X"e4061800",
		16#3959# => X"10000066",
		16#395a# => X"b9080082",
		16#395b# => X"84e60004",
		16#395c# => X"9d00fffc",
		16#395d# => X"e0e74003",
		16#395e# => X"e4853800",
		16#395f# => X"10000009",
		16#3960# => X"15000000",
		16#3961# => X"0000000c",
		16#3962# => X"8466000c",
		16#3963# => X"84e60004",
		16#3964# => X"e0e75803",
		16#3965# => X"e4853800",
		16#3966# => X"0c000006",
		16#3967# => X"15000000",
		16#3968# => X"84c60008",
		16#3969# => X"e4033000",
		16#396a# => X"0ffffff9",
		16#396b# => X"9d60fffc",
		16#396c# => X"8466000c",
		16#396d# => X"d404180c",
		16#396e# => X"d4043008",
		16#396f# => X"d4032008",
		16#3970# => X"d406200c",
		16#3971# => X"9c21000c",
		16#3972# => X"a8620000",
		16#3973# => X"8521fffc",
		16#3974# => X"8441fff4",
		16#3975# => X"03ffe737",
		16#3976# => X"85c1fff8",
		16#3977# => X"9c21000c",
		16#3978# => X"8521fffc",
		16#3979# => X"8441fff4",
		16#397a# => X"44004800",
		16#397b# => X"85c1fff8",
		16#397c# => X"19000001",
		16#397d# => X"84660008",
		16#397e# => X"a9086810",
		16#397f# => X"e4234000",
		16#3980# => X"13ffffc1",
		16#3981# => X"15000000",
		16#3982# => X"a8e50001",
		16#3983# => X"e0c42800",
		16#3984# => X"d403200c",
		16#3985# => X"d4032008",
		16#3986# => X"d404180c",
		16#3987# => X"d4041808",
		16#3988# => X"d4043804",
		16#3989# => X"03ffffe8",
		16#398a# => X"d4062800",
		16#398b# => X"b8a50043",
		16#398c# => X"19600001",
		16#398d# => X"b8650082",
		16#398e# => X"b8a50003",
		16#398f# => X"a96b6808",
		16#3990# => X"e0c61808",
		16#3991# => X"e0a55800",
		16#3992# => X"85070004",
		16#3993# => X"84650008",
		16#3994# => X"e0c83004",
		16#3995# => X"d4041808",
		16#3996# => X"d404280c",
		16#3997# => X"d403200c",
		16#3998# => X"d4073004",
		16#3999# => X"d4052008",
		16#399a# => X"9c21000c",
		16#399b# => X"a8620000",
		16#399c# => X"8521fffc",
		16#399d# => X"8441fff4",
		16#399e# => X"03ffe70e",
		16#399f# => X"85c1fff8",
		16#39a0# => X"a5080001",
		16#39a1# => X"bc280000",
		16#39a2# => X"10000009",
		16#39a3# => X"e0a32800",
		16#39a4# => X"84640000",
		16#39a5# => X"e0841802",
		16#39a6# => X"e0a51800",
		16#39a7# => X"84c40008",
		16#39a8# => X"8464000c",
		16#39a9# => X"d406180c",
		16#39aa# => X"d4033008",
		16#39ab# => X"a8650001",
		16#39ac# => X"d4072008",
		16#39ad# => X"d4041804",
		16#39ae# => X"18600001",
		16#39af# => X"a8636c10",
		16#39b0# => X"84630000",
		16#39b1# => X"e4851800",
		16#39b2# => X"13ffffbf",
		16#39b3# => X"18800001",
		16#39b4# => X"a8620000",
		16#39b5# => X"a8847a78",
		16#39b6# => X"07ffff09",
		16#39b7# => X"84840000",
		16#39b8# => X"03ffffba",
		16#39b9# => X"9c21000c",
		16#39ba# => X"1000000c",
		16#39bb# => X"bc430054",
		16#39bc# => X"9d03005b",
		16#39bd# => X"03ffff97",
		16#39be# => X"b8680003",
		16#39bf# => X"9c600001",
		16#39c0# => X"85670004",
		16#39c1# => X"e0a34008",
		16#39c2# => X"a8660000",
		16#39c3# => X"e0ab2804",
		16#39c4# => X"03ffffa9",
		16#39c5# => X"d4072804",
		16#39c6# => X"10000006",
		16#39c7# => X"bc430154",
		16#39c8# => X"b905004c",
		16#39c9# => X"9d08006e",
		16#39ca# => X"03ffff8a",
		16#39cb# => X"b8680003",
		16#39cc# => X"10000006",
		16#39cd# => X"bc430554",
		16#39ce# => X"b905004f",
		16#39cf# => X"9d080077",
		16#39d0# => X"03ffff84",
		16#39d1# => X"b8680003",
		16#39d2# => X"10000006",
		16#39d3# => X"15000000",
		16#39d4# => X"b9050052",
		16#39d5# => X"9d08007c",
		16#39d6# => X"03ffff7e",
		16#39d7# => X"b8680003",
		16#39d8# => X"9c6003f0",
		16#39d9# => X"03ffff7b",
		16#39da# => X"9d00007e",
		16#39db# => X"d7e117d4",
		16#39dc# => X"d7e197e0",
		16#39dd# => X"d7e1e7f4",
		16#39de# => X"d7e14ffc",
		16#39df# => X"d7e177d8",
		16#39e0# => X"d7e187dc",
		16#39e1# => X"d7e1a7e4",
		16#39e2# => X"d7e1b7e8",
		16#39e3# => X"d7e1c7ec",
		16#39e4# => X"d7e1d7f0",
		16#39e5# => X"d7e1f7f8",
		16#39e6# => X"85650008",
		16#39e7# => X"9c21ffd4",
		16#39e8# => X"aa450000",
		16#39e9# => X"ab830000",
		16#39ea# => X"bc0b0000",
		16#39eb# => X"10000027",
		16#39ec# => X"a8440000",
		16#39ed# => X"9864000c",
		16#39ee# => X"a483ffff",
		16#39ef# => X"a4a40008",
		16#39f0# => X"bc050000",
		16#39f1# => X"1000002e",
		16#39f2# => X"15000000",
		16#39f3# => X"84a20010",
		16#39f4# => X"bc250000",
		16#39f5# => X"0c00002a",
		16#39f6# => X"a4a40002",
		16#39f7# => X"bc050000",
		16#39f8# => X"10000033",
		16#39f9# => X"86120000",
		16#39fa# => X"9ec00000",
		16#39fb# => X"a9d60000",
		16#39fc# => X"a8b60000",
		16#39fd# => X"bc0e0000",
		16#39fe# => X"10000067",
		16#39ff# => X"a87c0000",
		16#3a00# => X"a8ce0000",
		16#3a01# => X"bcae0400",
		16#3a02# => X"10000003",
		16#3a03# => X"8482001c",
		16#3a04# => X"9cc00400",
		16#3a05# => X"85620024",
		16#3a06# => X"48005800",
		16#3a07# => X"15000000",
		16#3a08# => X"bdab0000",
		16#3a09# => X"100000c8",
		16#3a0a# => X"e2d65800",
		16#3a0b# => X"86920008",
		16#3a0c# => X"e2945802",
		16#3a0d# => X"e1ce5802",
		16#3a0e# => X"bc340000",
		16#3a0f# => X"13ffffed",
		16#3a10# => X"d412a008",
		16#3a11# => X"a9740000",
		16#3a12# => X"9c21002c",
		16#3a13# => X"8521fffc",
		16#3a14# => X"8441ffd4",
		16#3a15# => X"85c1ffd8",
		16#3a16# => X"8601ffdc",
		16#3a17# => X"8641ffe0",
		16#3a18# => X"8681ffe4",
		16#3a19# => X"86c1ffe8",
		16#3a1a# => X"8701ffec",
		16#3a1b# => X"8741fff0",
		16#3a1c# => X"8781fff4",
		16#3a1d# => X"44004800",
		16#3a1e# => X"87c1fff8",
		16#3a1f# => X"a87c0000",
		16#3a20# => X"07fff3c6",
		16#3a21# => X"a8820000",
		16#3a22# => X"bc2b0000",
		16#3a23# => X"10000122",
		16#3a24# => X"15000000",
		16#3a25# => X"9862000c",
		16#3a26# => X"a483ffff",
		16#3a27# => X"a4a40002",
		16#3a28# => X"bc050000",
		16#3a29# => X"0fffffd1",
		16#3a2a# => X"86120000",
		16#3a2b# => X"a6c40001",
		16#3a2c# => X"bc160000",
		16#3a2d# => X"1000003f",
		16#3a2e# => X"a9d60000",
		16#3a2f# => X"aac50000",
		16#3a30# => X"abc50000",
		16#3a31# => X"ab450000",
		16#3a32# => X"aa850000",
		16#3a33# => X"bc140000",
		16#3a34# => X"1000002c",
		16#3a35# => X"bc3e0000",
		16#3a36# => X"0c000102",
		16#3a37# => X"a87a0000",
		16#3a38# => X"e4b6a000",
		16#3a39# => X"10000003",
		16#3a3a# => X"ab160000",
		16#3a3b# => X"ab140000",
		16#3a3c# => X"84c20014",
		16#3a3d# => X"85c20008",
		16#3a3e# => X"84620000",
		16#3a3f# => X"e1c67000",
		16#3a40# => X"e5587000",
		16#3a41# => X"10000003",
		16#3a42# => X"9c800001",
		16#3a43# => X"9c800000",
		16#3a44# => X"a48400ff",
		16#3a45# => X"bc040000",
		16#3a46# => X"0c0000db",
		16#3a47# => X"e5983000",
		16#3a48# => X"100000c5",
		16#3a49# => X"a89a0000",
		16#3a4a# => X"85620024",
		16#3a4b# => X"a87c0000",
		16#3a4c# => X"8482001c",
		16#3a4d# => X"48005800",
		16#3a4e# => X"a8ba0000",
		16#3a4f# => X"bdab0000",
		16#3a50# => X"10000081",
		16#3a51# => X"a9cb0000",
		16#3a52# => X"e2d67002",
		16#3a53# => X"bc360000",
		16#3a54# => X"0c0000c6",
		16#3a55# => X"a87c0000",
		16#3a56# => X"85720008",
		16#3a57# => X"e35a7000",
		16#3a58# => X"e16b7002",
		16#3a59# => X"e2947002",
		16#3a5a# => X"bc2b0000",
		16#3a5b# => X"0fffffb7",
		16#3a5c# => X"d4125808",
		16#3a5d# => X"bc140000",
		16#3a5e# => X"0fffffd8",
		16#3a5f# => X"bc3e0000",
		16#3a60# => X"87500000",
		16#3a61# => X"86900004",
		16#3a62# => X"9fc00000",
		16#3a63# => X"03ffffd0",
		16#3a64# => X"9e100008",
		16#3a65# => X"86d00000",
		16#3a66# => X"85d00004",
		16#3a67# => X"03ffff95",
		16#3a68# => X"9e100008",
		16#3a69# => X"86d00000",
		16#3a6a# => X"85d00004",
		16#3a6b# => X"9e100008",
		16#3a6c# => X"bc0e0000",
		16#3a6d# => X"13fffffc",
		16#3a6e# => X"15000000",
		16#3a6f# => X"a463ffff",
		16#3a70# => X"a4830200",
		16#3a71# => X"bc040000",
		16#3a72# => X"10000023",
		16#3a73# => X"86820008",
		16#3a74# => X"e48ea000",
		16#3a75# => X"10000038",
		16#3a76# => X"ab540000",
		16#3a77# => X"a4830480",
		16#3a78# => X"bc240000",
		16#3a79# => X"1000005d",
		16#3a7a# => X"abd40000",
		16#3a7b# => X"84620000",
		16#3a7c# => X"aa8e0000",
		16#3a7d# => X"a8960000",
		16#3a7e# => X"a8ba0000",
		16#3a7f# => X"0400027b",
		16#3a80# => X"ab0e0000",
		16#3a81# => X"84820008",
		16#3a82# => X"84620000",
		16#3a83# => X"e3c4f002",
		16#3a84# => X"e343d000",
		16#3a85# => X"d402f008",
		16#3a86# => X"d402d000",
		16#3a87# => X"84720008",
		16#3a88# => X"e2d6c000",
		16#3a89# => X"e283a002",
		16#3a8a# => X"e1cec002",
		16#3a8b# => X"bc340000",
		16#3a8c# => X"0fffff85",
		16#3a8d# => X"d412a008",
		16#3a8e# => X"bc0e0000",
		16#3a8f# => X"0fffffe0",
		16#3a90# => X"9862000c",
		16#3a91# => X"86d00000",
		16#3a92# => X"85d00004",
		16#3a93# => X"03ffffd9",
		16#3a94# => X"9e100008",
		16#3a95# => X"84620000",
		16#3a96# => X"ab140000",
		16#3a97# => X"e4947000",
		16#3a98# => X"10000003",
		16#3a99# => X"9ca00001",
		16#3a9a# => X"a8a40000",
		16#3a9b# => X"a4a500ff",
		16#3a9c# => X"bc050000",
		16#3a9d# => X"0c000020",
		16#3a9e# => X"15000000",
		16#3a9f# => X"84c20014",
		16#3aa0# => X"e48e3000",
		16#3aa1# => X"10000011",
		16#3aa2# => X"a8960000",
		16#3aa3# => X"85620024",
		16#3aa4# => X"a87c0000",
		16#3aa5# => X"8482001c",
		16#3aa6# => X"48005800",
		16#3aa7# => X"a8b60000",
		16#3aa8# => X"bdab0000",
		16#3aa9# => X"10000028",
		16#3aaa# => X"aa8b0000",
		16#3aab# => X"03ffffdc",
		16#3aac# => X"ab0b0000",
		16#3aad# => X"abce0000",
		16#3aae# => X"84620000",
		16#3aaf# => X"ab4e0000",
		16#3ab0# => X"03ffffcd",
		16#3ab1# => X"aa8e0000",
		16#3ab2# => X"a8ae0000",
		16#3ab3# => X"04000247",
		16#3ab4# => X"aa8e0000",
		16#3ab5# => X"84820008",
		16#3ab6# => X"84620000",
		16#3ab7# => X"e0847002",
		16#3ab8# => X"e0637000",
		16#3ab9# => X"d4022008",
		16#3aba# => X"d4021800",
		16#3abb# => X"03ffffcc",
		16#3abc# => X"ab0e0000",
		16#3abd# => X"84a20010",
		16#3abe# => X"e4432800",
		16#3abf# => X"10000003",
		16#3ac0# => X"9c800001",
		16#3ac1# => X"9c800000",
		16#3ac2# => X"a48400ff",
		16#3ac3# => X"bc040000",
		16#3ac4# => X"13ffffdb",
		16#3ac5# => X"a8960000",
		16#3ac6# => X"04000234",
		16#3ac7# => X"a8b40000",
		16#3ac8# => X"84a20000",
		16#3ac9# => X"a87c0000",
		16#3aca# => X"e0a5a000",
		16#3acb# => X"a8820000",
		16#3acc# => X"07fffc14",
		16#3acd# => X"d4022800",
		16#3ace# => X"bc2b0000",
		16#3acf# => X"0fffffb8",
		16#3ad0# => X"15000000",
		16#3ad1# => X"9462000c",
		16#3ad2# => X"a8630040",
		16#3ad3# => X"9d60ffff",
		16#3ad4# => X"03ffff3e",
		16#3ad5# => X"dc02180c",
		16#3ad6# => X"84a20014",
		16#3ad7# => X"84820010",
		16#3ad8# => X"e0c52800",
		16#3ad9# => X"87420000",
		16#3ada# => X"e0a62800",
		16#3adb# => X"e35a2002",
		16#3adc# => X"ba85005f",
		16#3add# => X"9cda0001",
		16#3ade# => X"e0b42800",
		16#3adf# => X"e0c67000",
		16#3ae0# => X"ba850081",
		16#3ae1# => X"e4743000",
		16#3ae2# => X"10000004",
		16#3ae3# => X"a8b40000",
		16#3ae4# => X"aa860000",
		16#3ae5# => X"a8a60000",
		16#3ae6# => X"a4630400",
		16#3ae7# => X"bc030000",
		16#3ae8# => X"1000001a",
		16#3ae9# => X"a87c0000",
		16#3aea# => X"07ffe370",
		16#3aeb# => X"a8850000",
		16#3aec# => X"bc2b0000",
		16#3aed# => X"0c00001d",
		16#3aee# => X"ab0b0000",
		16#3aef# => X"a86b0000",
		16#3af0# => X"84820010",
		16#3af1# => X"040001c5",
		16#3af2# => X"a8ba0000",
		16#3af3# => X"9462000c",
		16#3af4# => X"9c80fb7f",
		16#3af5# => X"e0632003",
		16#3af6# => X"a8630080",
		16#3af7# => X"dc02180c",
		16#3af8# => X"e078d000",
		16#3af9# => X"e354d002",
		16#3afa# => X"d402a014",
		16#3afb# => X"d402d008",
		16#3afc# => X"d402c010",
		16#3afd# => X"d4021800",
		16#3afe# => X"abce0000",
		16#3aff# => X"ab4e0000",
		16#3b00# => X"03ffff7d",
		16#3b01# => X"aa8e0000",
		16#3b02# => X"04000736",
		16#3b03# => X"a87c0000",
		16#3b04# => X"bc2b0000",
		16#3b05# => X"13fffff3",
		16#3b06# => X"ab0b0000",
		16#3b07# => X"a87c0000",
		16#3b08# => X"07fffe07",
		16#3b09# => X"84820010",
		16#3b0a# => X"9c60000c",
		16#3b0b# => X"03ffffc6",
		16#3b0c# => X"d41c1800",
		16#3b0d# => X"a8b80000",
		16#3b0e# => X"040001ec",
		16#3b0f# => X"a9d80000",
		16#3b10# => X"84620008",
		16#3b11# => X"84820000",
		16#3b12# => X"e063c002",
		16#3b13# => X"e304c000",
		16#3b14# => X"e2d67002",
		16#3b15# => X"d4021808",
		16#3b16# => X"bc360000",
		16#3b17# => X"13ffff3f",
		16#3b18# => X"d402c000",
		16#3b19# => X"a87c0000",
		16#3b1a# => X"07fffbc6",
		16#3b1b# => X"a8820000",
		16#3b1c# => X"bc2b0000",
		16#3b1d# => X"13ffffb4",
		16#3b1e# => X"15000000",
		16#3b1f# => X"03ffff37",
		16#3b20# => X"abd60000",
		16#3b21# => X"84a20010",
		16#3b22# => X"e4432800",
		16#3b23# => X"10000003",
		16#3b24# => X"9c800001",
		16#3b25# => X"9c800000",
		16#3b26# => X"a48400ff",
		16#3b27# => X"bc040000",
		16#3b28# => X"13ffff20",
		16#3b29# => X"e5983000",
		16#3b2a# => X"a89a0000",
		16#3b2b# => X"040001cf",
		16#3b2c# => X"a8ae0000",
		16#3b2d# => X"84a20000",
		16#3b2e# => X"a87c0000",
		16#3b2f# => X"e0a57000",
		16#3b30# => X"a8820000",
		16#3b31# => X"07fffbaf",
		16#3b32# => X"d4022800",
		16#3b33# => X"bc2b0000",
		16#3b34# => X"0fffff1f",
		16#3b35# => X"e2d67002",
		16#3b36# => X"03ffff9c",
		16#3b37# => X"9462000c",
		16#3b38# => X"9c80000a",
		16#3b39# => X"04000132",
		16#3b3a# => X"a8b40000",
		16#3b3b# => X"bc0b0000",
		16#3b3c# => X"10000006",
		16#3b3d# => X"15000000",
		16#3b3e# => X"9ecb0001",
		16#3b3f# => X"9fc00001",
		16#3b40# => X"03fffef8",
		16#3b41# => X"e2d6d002",
		16#3b42# => X"9ed40001",
		16#3b43# => X"03fffef5",
		16#3b44# => X"9fc00001",
		16#3b45# => X"9462000c",
		16#3b46# => X"a8630040",
		16#3b47# => X"9d60ffff",
		16#3b48# => X"dc02180c",
		16#3b49# => X"9c400009",
		16#3b4a# => X"03fffec8",
		16#3b4b# => X"d41c1000",
		16#3b4c# => X"d7e187f0",
		16#3b4d# => X"d7e197f4",
		16#3b4e# => X"d7e1a7f8",
		16#3b4f# => X"d7e14ffc",
		16#3b50# => X"d7e117e8",
		16#3b51# => X"d7e177ec",
		16#3b52# => X"9c21ffe8",
		16#3b53# => X"9e0302e0",
		16#3b54# => X"07fffd4f",
		16#3b55# => X"aa840000",
		16#3b56# => X"bc100000",
		16#3b57# => X"1000001c",
		16#3b58# => X"aa500000",
		16#3b59# => X"9e400000",
		16#3b5a# => X"85d00004",
		16#3b5b# => X"9dceffff",
		16#3b5c# => X"bd8e0000",
		16#3b5d# => X"10000012",
		16#3b5e# => X"84500008",
		16#3b5f# => X"9c42000c",
		16#3b60# => X"98620000",
		16#3b61# => X"9dceffff",
		16#3b62# => X"bc030000",
		16#3b63# => X"10000009",
		16#3b64# => X"9c62fff4",
		16#3b65# => X"98a20002",
		16#3b66# => X"bc05ffff",
		16#3b67# => X"10000006",
		16#3b68# => X"bd6e0000",
		16#3b69# => X"4800a000",
		16#3b6a# => X"15000000",
		16#3b6b# => X"e2525804",
		16#3b6c# => X"bd6e0000",
		16#3b6d# => X"13fffff3",
		16#3b6e# => X"9c420068",
		16#3b6f# => X"86100000",
		16#3b70# => X"bc300000",
		16#3b71# => X"13ffffe9",
		16#3b72# => X"15000000",
		16#3b73# => X"07fffd32",
		16#3b74# => X"15000000",
		16#3b75# => X"9c210018",
		16#3b76# => X"a9720000",
		16#3b77# => X"8521fffc",
		16#3b78# => X"8441ffe8",
		16#3b79# => X"85c1ffec",
		16#3b7a# => X"8601fff0",
		16#3b7b# => X"8641fff4",
		16#3b7c# => X"44004800",
		16#3b7d# => X"8681fff8",
		16#3b7e# => X"d7e187ec",
		16#3b7f# => X"d7e197f0",
		16#3b80# => X"d7e1a7f4",
		16#3b81# => X"d7e1b7f8",
		16#3b82# => X"d7e14ffc",
		16#3b83# => X"d7e117e4",
		16#3b84# => X"d7e177e8",
		16#3b85# => X"9c21ffe4",
		16#3b86# => X"9e0302e0",
		16#3b87# => X"aa830000",
		16#3b88# => X"07fffd1b",
		16#3b89# => X"aac40000",
		16#3b8a# => X"bc100000",
		16#3b8b# => X"1000001c",
		16#3b8c# => X"aa500000",
		16#3b8d# => X"9e400000",
		16#3b8e# => X"85d00004",
		16#3b8f# => X"9dceffff",
		16#3b90# => X"bd8e0000",
		16#3b91# => X"10000012",
		16#3b92# => X"84500008",
		16#3b93# => X"9c42000c",
		16#3b94# => X"98a20000",
		16#3b95# => X"9dceffff",
		16#3b96# => X"bc050000",
		16#3b97# => X"10000009",
		16#3b98# => X"9c82fff4",
		16#3b99# => X"98a20002",
		16#3b9a# => X"bc05ffff",
		16#3b9b# => X"10000005",
		16#3b9c# => X"a8740000",
		16#3b9d# => X"4800b000",
		16#3b9e# => X"15000000",
		16#3b9f# => X"e2525804",
		16#3ba0# => X"bd6e0000",
		16#3ba1# => X"13fffff3",
		16#3ba2# => X"9c420068",
		16#3ba3# => X"86100000",
		16#3ba4# => X"bc300000",
		16#3ba5# => X"13ffffe9",
		16#3ba6# => X"15000000",
		16#3ba7# => X"07fffcfe",
		16#3ba8# => X"15000000",
		16#3ba9# => X"9c21001c",
		16#3baa# => X"a9720000",
		16#3bab# => X"8521fffc",
		16#3bac# => X"8441ffe4",
		16#3bad# => X"85c1ffe8",
		16#3bae# => X"8601ffec",
		16#3baf# => X"8641fff0",
		16#3bb0# => X"8681fff4",
		16#3bb1# => X"44004800",
		16#3bb2# => X"86c1fff8",
		16#3bb3# => X"d7e117f4",
		16#3bb4# => X"d7e177f8",
		16#3bb5# => X"d7e14ffc",
		16#3bb6# => X"19c00001",
		16#3bb7# => X"9c21fff4",
		16#3bb8# => X"a8450000",
		16#3bb9# => X"bc050000",
		16#3bba# => X"10000009",
		16#3bbb# => X"a9ce3ea4",
		16#3bbc# => X"18800001",
		16#3bbd# => X"a8650000",
		16#3bbe# => X"04000972",
		16#3bbf# => X"a88440d0",
		16#3bc0# => X"bc0b0000",
		16#3bc1# => X"0c000008",
		16#3bc2# => X"a8620000",
		16#3bc3# => X"9c21000c",
		16#3bc4# => X"a96e0000",
		16#3bc5# => X"8521fffc",
		16#3bc6# => X"8441fff4",
		16#3bc7# => X"44004800",
		16#3bc8# => X"85c1fff8",
		16#3bc9# => X"04000967",
		16#3bca# => X"a88e0000",
		16#3bcb# => X"bc0b0000",
		16#3bcc# => X"13fffff7",
		16#3bcd# => X"a8620000",
		16#3bce# => X"18800001",
		16#3bcf# => X"a8843b54",
		16#3bd0# => X"04000960",
		16#3bd1# => X"9dc00000",
		16#3bd2# => X"e42b7000",
		16#3bd3# => X"13fffff0",
		16#3bd4# => X"15000000",
		16#3bd5# => X"19c00001",
		16#3bd6# => X"03ffffed",
		16#3bd7# => X"a9ce3ea4",
		16#3bd8# => X"19600001",
		16#3bd9# => X"44004800",
		16#3bda# => X"a96b6db4",
		16#3bdb# => X"19600001",
		16#3bdc# => X"44004800",
		16#3bdd# => X"a96b6d94",
		16#3bde# => X"44004800",
		16#3bdf# => X"9d600000",
		16#3be0# => X"19600001",
		16#3be1# => X"44004800",
		16#3be2# => X"a96b40d8",
		16#3be3# => X"a8a40000",
		16#3be4# => X"a8830000",
		16#3be5# => X"18600001",
		16#3be6# => X"d7e14ffc",
		16#3be7# => X"a86363e0",
		16#3be8# => X"9c21fffc",
		16#3be9# => X"84630000",
		16#3bea# => X"9c210004",
		16#3beb# => X"8521fffc",
		16#3bec# => X"03ffffc7",
		16#3bed# => X"15000000",
		16#3bee# => X"19600001",
		16#3bef# => X"44004800",
		16#3bf0# => X"a96b40d8",
		16#3bf1# => X"98a4000c",
		16#3bf2# => X"a4c5ffff",
		16#3bf3# => X"d7e117ec",
		16#3bf4# => X"d7e177f0",
		16#3bf5# => X"d7e14ffc",
		16#3bf6# => X"d7e187f4",
		16#3bf7# => X"d7e197f8",
		16#3bf8# => X"a8440000",
		16#3bf9# => X"a4860002",
		16#3bfa# => X"9c21ffb0",
		16#3bfb# => X"bc040000",
		16#3bfc# => X"0c000039",
		16#3bfd# => X"a9c30000",
		16#3bfe# => X"9882000e",
		16#3bff# => X"bd840000",
		16#3c00# => X"10000018",
		16#3c01# => X"a4c60080",
		16#3c02# => X"04000f0e",
		16#3c03# => X"a8a10000",
		16#3c04# => X"bd6b0000",
		16#3c05# => X"0c000010",
		16#3c06# => X"84810004",
		16#3c07# => X"a8a08000",
		16#3c08# => X"a484f000",
		16#3c09# => X"ac642000",
		16#3c0a# => X"e4242800",
		16#3c0b# => X"e2401802",
		16#3c0c# => X"e2521804",
		16#3c0d# => X"ae52ffff",
		16#3c0e# => X"0c000045",
		16#3c0f# => X"ba52005f",
		16#3c10# => X"9462000c",
		16#3c11# => X"a8630800",
		16#3c12# => X"9e000400",
		16#3c13# => X"0000000b",
		16#3c14# => X"dc02180c",
		16#3c15# => X"98a2000c",
		16#3c16# => X"a4c5ffff",
		16#3c17# => X"a4c60080",
		16#3c18# => X"bc260000",
		16#3c19# => X"0c000038",
		16#3c1a# => X"9e000040",
		16#3c1b# => X"a8a50800",
		16#3c1c# => X"9e400000",
		16#3c1d# => X"dc02280c",
		16#3c1e# => X"a86e0000",
		16#3c1f# => X"07ffe23b",
		16#3c20# => X"a8900000",
		16#3c21# => X"bc2b0000",
		16#3c22# => X"0c00003d",
		16#3c23# => X"18800000",
		16#3c24# => X"9462000c",
		16#3c25# => X"a8630080",
		16#3c26# => X"a884df10",
		16#3c27# => X"bc120000",
		16#3c28# => X"d40e203c",
		16#3c29# => X"dc02180c",
		16#3c2a# => X"d4025800",
		16#3c2b# => X"d4025810",
		16#3c2c# => X"0c000015",
		16#3c2d# => X"d4028014",
		16#3c2e# => X"9c210050",
		16#3c2f# => X"8521fffc",
		16#3c30# => X"8441ffec",
		16#3c31# => X"85c1fff0",
		16#3c32# => X"8601fff4",
		16#3c33# => X"44004800",
		16#3c34# => X"8641fff8",
		16#3c35# => X"9c620043",
		16#3c36# => X"d4021800",
		16#3c37# => X"d4021810",
		16#3c38# => X"9c600001",
		16#3c39# => X"d4021814",
		16#3c3a# => X"9c210050",
		16#3c3b# => X"8521fffc",
		16#3c3c# => X"8441ffec",
		16#3c3d# => X"85c1fff0",
		16#3c3e# => X"8601fff4",
		16#3c3f# => X"44004800",
		16#3c40# => X"8641fff8",
		16#3c41# => X"9882000e",
		16#3c42# => X"04000eec",
		16#3c43# => X"a86e0000",
		16#3c44# => X"bc0b0000",
		16#3c45# => X"13ffffe9",
		16#3c46# => X"15000000",
		16#3c47# => X"9462000c",
		16#3c48# => X"a8630001",
		16#3c49# => X"dc02180c",
		16#3c4a# => X"9c210050",
		16#3c4b# => X"8521fffc",
		16#3c4c# => X"8441ffec",
		16#3c4d# => X"85c1fff0",
		16#3c4e# => X"8601fff4",
		16#3c4f# => X"44004800",
		16#3c50# => X"8641fff8",
		16#3c51# => X"03ffffca",
		16#3c52# => X"9e000400",
		16#3c53# => X"18800001",
		16#3c54# => X"84620028",
		16#3c55# => X"a8841444",
		16#3c56# => X"e4232000",
		16#3c57# => X"13ffffb9",
		16#3c58# => X"15000000",
		16#3c59# => X"9462000c",
		16#3c5a# => X"9e000400",
		16#3c5b# => X"e0638004",
		16#3c5c# => X"d402804c",
		16#3c5d# => X"03ffffc1",
		16#3c5e# => X"dc02180c",
		16#3c5f# => X"9862000c",
		16#3c60# => X"a4830200",
		16#3c61# => X"bc240000",
		16#3c62# => X"13ffffcc",
		16#3c63# => X"a8630002",
		16#3c64# => X"9c820043",
		16#3c65# => X"dc02180c",
		16#3c66# => X"9c600001",
		16#3c67# => X"d4022000",
		16#3c68# => X"d4022010",
		16#3c69# => X"03ffffc5",
		16#3c6a# => X"d4021814",
		16#3c6b# => X"d7e117fc",
		16#3c6c# => X"a4c30003",
		16#3c6d# => X"9c21fffc",
		16#3c6e# => X"bc060000",
		16#3c6f# => X"10000016",
		16#3c70# => X"a48400ff",
		16#3c71# => X"bc050000",
		16#3c72# => X"10000027",
		16#3c73# => X"a9650000",
		16#3c74# => X"8cc30000",
		16#3c75# => X"e4062000",
		16#3c76# => X"10000023",
		16#3c77# => X"a9630000",
		16#3c78# => X"00000008",
		16#3c79# => X"9ca5ffff",
		16#3c7a# => X"1000001f",
		16#3c7b# => X"a9650000",
		16#3c7c# => X"8cc30000",
		16#3c7d# => X"e4062000",
		16#3c7e# => X"1000001e",
		16#3c7f# => X"9ca5ffff",
		16#3c80# => X"9c630001",
		16#3c81# => X"a4c30003",
		16#3c82# => X"bc260000",
		16#3c83# => X"13fffff7",
		16#3c84# => X"bc050000",
		16#3c85# => X"bca50003",
		16#3c86# => X"0c00001a",
		16#3c87# => X"b8c40008",
		16#3c88# => X"bc050000",
		16#3c89# => X"10000010",
		16#3c8a# => X"a9650000",
		16#3c8b# => X"8cc30000",
		16#3c8c# => X"e4062000",
		16#3c8d# => X"1000000c",
		16#3c8e# => X"a9630000",
		16#3c8f# => X"00000006",
		16#3c90# => X"9ca5ffff",
		16#3c91# => X"8cc30000",
		16#3c92# => X"e4062000",
		16#3c93# => X"10000009",
		16#3c94# => X"9ca5ffff",
		16#3c95# => X"bc250000",
		16#3c96# => X"13fffffb",
		16#3c97# => X"9c630001",
		16#3c98# => X"a9650000",
		16#3c99# => X"9c210004",
		16#3c9a# => X"44004800",
		16#3c9b# => X"8441fffc",
		16#3c9c# => X"9c210004",
		16#3c9d# => X"a9630000",
		16#3c9e# => X"44004800",
		16#3c9f# => X"8441fffc",
		16#3ca0# => X"e0c62004",
		16#3ca1# => X"b9060010",
		16#3ca2# => X"e1083004",
		16#3ca3# => X"84c30000",
		16#3ca4# => X"1840fefe",
		16#3ca5# => X"e0c83005",
		16#3ca6# => X"a842feff",
		16#3ca7# => X"e0e61000",
		16#3ca8# => X"acc6ffff",
		16#3ca9# => X"18408080",
		16#3caa# => X"e0c73003",
		16#3cab# => X"a8428080",
		16#3cac# => X"e0c61003",
		16#3cad# => X"bc260000",
		16#3cae# => X"13ffffdb",
		16#3caf# => X"bc050000",
		16#3cb0# => X"9ca5fffc",
		16#3cb1# => X"bc450003",
		16#3cb2# => X"13fffff1",
		16#3cb3# => X"9c630004",
		16#3cb4# => X"03ffffd5",
		16#3cb5# => X"bc050000",
		16#3cb6# => X"a9030000",
		16#3cb7# => X"a9840000",
		16#3cb8# => X"bca5000f",
		16#3cb9# => X"10000007",
		16#3cba# => X"a8e50000",
		16#3cbb# => X"e0c41804",
		16#3cbc# => X"a4c60003",
		16#3cbd# => X"bc260000",
		16#3cbe# => X"0c00000f",
		16#3cbf# => X"a8c40000",
		16#3cc0# => X"bc070000",
		16#3cc1# => X"1000000a",
		16#3cc2# => X"15000000",
		16#3cc3# => X"9c800000",
		16#3cc4# => X"e0cc2000",
		16#3cc5# => X"e0a82000",
		16#3cc6# => X"8cc60000",
		16#3cc7# => X"9c840001",
		16#3cc8# => X"e4243800",
		16#3cc9# => X"13fffffb",
		16#3cca# => X"d8053000",
		16#3ccb# => X"44004800",
		16#3ccc# => X"a9630000",
		16#3ccd# => X"a9050000",
		16#3cce# => X"a8e30000",
		16#3ccf# => X"85660000",
		16#3cd0# => X"9d08fff0",
		16#3cd1# => X"d4075800",
		16#3cd2# => X"bc48000f",
		16#3cd3# => X"85660004",
		16#3cd4# => X"d4075804",
		16#3cd5# => X"85660008",
		16#3cd6# => X"d4075808",
		16#3cd7# => X"8566000c",
		16#3cd8# => X"9cc60010",
		16#3cd9# => X"d407580c",
		16#3cda# => X"13fffff5",
		16#3cdb# => X"9ce70010",
		16#3cdc# => X"9ca5fff0",
		16#3cdd# => X"b8c50044",
		16#3cde# => X"9d860001",
		16#3cdf# => X"b8c60004",
		16#3ce0# => X"b98c0004",
		16#3ce1# => X"e0a53002",
		16#3ce2# => X"e1036000",
		16#3ce3# => X"a8e50000",
		16#3ce4# => X"bca50003",
		16#3ce5# => X"13ffffdb",
		16#3ce6# => X"e1846000",
		16#3ce7# => X"9c800000",
		16#3ce8# => X"e0cc2000",
		16#3ce9# => X"e0e82000",
		16#3cea# => X"84c60000",
		16#3ceb# => X"9c840004",
		16#3cec# => X"d4073000",
		16#3ced# => X"e0c52002",
		16#3cee# => X"bc460003",
		16#3cef# => X"13fffffa",
		16#3cf0# => X"e0cc2000",
		16#3cf1# => X"9ca5fffc",
		16#3cf2# => X"b8e50042",
		16#3cf3# => X"9c870001",
		16#3cf4# => X"b8e70002",
		16#3cf5# => X"b8840002",
		16#3cf6# => X"e0e53802",
		16#3cf7# => X"e1082000",
		16#3cf8# => X"03ffffc8",
		16#3cf9# => X"e18c2000",
		16#3cfa# => X"d7e117fc",
		16#3cfb# => X"a9030000",
		16#3cfc# => X"9c21fffc",
		16#3cfd# => X"a9640000",
		16#3cfe# => X"e4a32000",
		16#3cff# => X"10000016",
		16#3d00# => X"a8e50000",
		16#3d01# => X"e0c42800",
		16#3d02# => X"e4633000",
		16#3d03# => X"10000013",
		16#3d04# => X"bca5000f",
		16#3d05# => X"bc050000",
		16#3d06# => X"1000000b",
		16#3d07# => X"15000000",
		16#3d08# => X"e0832800",
		16#3d09# => X"9ca5ffff",
		16#3d0a# => X"9cc6ffff",
		16#3d0b# => X"9c84ffff",
		16#3d0c# => X"8c460000",
		16#3d0d# => X"9ca5ffff",
		16#3d0e# => X"bc25ffff",
		16#3d0f# => X"13fffffb",
		16#3d10# => X"d8041000",
		16#3d11# => X"9c210004",
		16#3d12# => X"a9630000",
		16#3d13# => X"44004800",
		16#3d14# => X"8441fffc",
		16#3d15# => X"bca5000f",
		16#3d16# => X"0c000011",
		16#3d17# => X"e0c41804",
		16#3d18# => X"bc070000",
		16#3d19# => X"13fffff8",
		16#3d1a# => X"15000000",
		16#3d1b# => X"9c800000",
		16#3d1c# => X"e0cb2000",
		16#3d1d# => X"e0a82000",
		16#3d1e# => X"8cc60000",
		16#3d1f# => X"9c840001",
		16#3d20# => X"e4243800",
		16#3d21# => X"13fffffb",
		16#3d22# => X"d8053000",
		16#3d23# => X"9c210004",
		16#3d24# => X"a9630000",
		16#3d25# => X"44004800",
		16#3d26# => X"8441fffc",
		16#3d27# => X"a4c60003",
		16#3d28# => X"bc260000",
		16#3d29# => X"13fffff0",
		16#3d2a# => X"bc070000",
		16#3d2b# => X"a9050000",
		16#3d2c# => X"a8c40000",
		16#3d2d# => X"a8e30000",
		16#3d2e# => X"85660000",
		16#3d2f# => X"9d08fff0",
		16#3d30# => X"d4075800",
		16#3d31# => X"bc48000f",
		16#3d32# => X"85660004",
		16#3d33# => X"d4075804",
		16#3d34# => X"85660008",
		16#3d35# => X"d4075808",
		16#3d36# => X"8566000c",
		16#3d37# => X"9cc60010",
		16#3d38# => X"d407580c",
		16#3d39# => X"13fffff5",
		16#3d3a# => X"9ce70010",
		16#3d3b# => X"9ca5fff0",
		16#3d3c# => X"b8c50044",
		16#3d3d# => X"9d660001",
		16#3d3e# => X"b8c60004",
		16#3d3f# => X"b96b0004",
		16#3d40# => X"e0a53002",
		16#3d41# => X"e1035800",
		16#3d42# => X"a8e50000",
		16#3d43# => X"bca50003",
		16#3d44# => X"13ffffd4",
		16#3d45# => X"e1645800",
		16#3d46# => X"9c800000",
		16#3d47# => X"e0cb2000",
		16#3d48# => X"e0e82000",
		16#3d49# => X"84c60000",
		16#3d4a# => X"9c840004",
		16#3d4b# => X"d4073000",
		16#3d4c# => X"e0c52002",
		16#3d4d# => X"bc460003",
		16#3d4e# => X"13fffffa",
		16#3d4f# => X"e0cb2000",
		16#3d50# => X"9ca5fffc",
		16#3d51# => X"b8e50042",
		16#3d52# => X"9c870001",
		16#3d53# => X"b8e70002",
		16#3d54# => X"b8840002",
		16#3d55# => X"e0e53802",
		16#3d56# => X"e1082000",
		16#3d57# => X"03ffffc1",
		16#3d58# => X"e16b2000",
		16#3d59# => X"d7e117fc",
		16#3d5a# => X"a4e30003",
		16#3d5b# => X"9c21fffc",
		16#3d5c# => X"bc070000",
		16#3d5d# => X"10000011",
		16#3d5e# => X"a8c30000",
		16#3d5f# => X"bc050000",
		16#3d60# => X"10000045",
		16#3d61# => X"15000000",
		16#3d62# => X"b9040018",
		16#3d63# => X"9ca5ffff",
		16#3d64# => X"00000004",
		16#3d65# => X"b9080098",
		16#3d66# => X"1000003f",
		16#3d67# => X"9ca5ffff",
		16#3d68# => X"d8064000",
		16#3d69# => X"9cc60001",
		16#3d6a# => X"a4e60003",
		16#3d6b# => X"bc270000",
		16#3d6c# => X"13fffffa",
		16#3d6d# => X"bc050000",
		16#3d6e# => X"bca50003",
		16#3d6f# => X"1000002c",
		16#3d70# => X"bc050000",
		16#3d71# => X"a50400ff",
		16#3d72# => X"a8e60000",
		16#3d73# => X"b9680008",
		16#3d74# => X"bc45000f",
		16#3d75# => X"e10b4004",
		16#3d76# => X"b9680010",
		16#3d77# => X"0c000014",
		16#3d78# => X"e10b4004",
		16#3d79# => X"a8e60000",
		16#3d7a# => X"a9850000",
		16#3d7b# => X"d4074000",
		16#3d7c# => X"d4074004",
		16#3d7d# => X"d4074008",
		16#3d7e# => X"d407400c",
		16#3d7f# => X"9d8cfff0",
		16#3d80# => X"bc4c000f",
		16#3d81# => X"13fffffa",
		16#3d82# => X"9ce70010",
		16#3d83# => X"9ca5fff0",
		16#3d84# => X"9c40fff0",
		16#3d85# => X"e0e51003",
		16#3d86# => X"a4a5000f",
		16#3d87# => X"9ce70010",
		16#3d88# => X"bc450003",
		16#3d89# => X"0c000010",
		16#3d8a# => X"e0e63800",
		16#3d8b# => X"9cc00000",
		16#3d8c# => X"e1673000",
		16#3d8d# => X"9cc60004",
		16#3d8e# => X"d40b4000",
		16#3d8f# => X"e1653002",
		16#3d90# => X"bc4b0003",
		16#3d91# => X"13fffffc",
		16#3d92# => X"e1673000",
		16#3d93# => X"9ca5fffc",
		16#3d94# => X"9c40fffc",
		16#3d95# => X"e0c51003",
		16#3d96# => X"a4a50003",
		16#3d97# => X"9cc60004",
		16#3d98# => X"e0e73000",
		16#3d99# => X"a8c70000",
		16#3d9a# => X"bc050000",
		16#3d9b# => X"1000000a",
		16#3d9c# => X"15000000",
		16#3d9d# => X"b8840018",
		16#3d9e# => X"9ce00000",
		16#3d9f# => X"b9040098",
		16#3da0# => X"e0863800",
		16#3da1# => X"9ce70001",
		16#3da2# => X"e4253800",
		16#3da3# => X"13fffffd",
		16#3da4# => X"d8044000",
		16#3da5# => X"9c210004",
		16#3da6# => X"a9630000",
		16#3da7# => X"44004800",
		16#3da8# => X"8441fffc",
		16#3da9# => X"d7e117f4",
		16#3daa# => X"d7e177f8",
		16#3dab# => X"d7e14ffc",
		16#3dac# => X"a8440000",
		16#3dad# => X"8483004c",
		16#3dae# => X"9c21fff4",
		16#3daf# => X"bc240000",
		16#3db0# => X"0c000012",
		16#3db1# => X"a9c30000",
		16#3db2# => X"b8620002",
		16#3db3# => X"e0841800",
		16#3db4# => X"85640000",
		16#3db5# => X"bc0b0000",
		16#3db6# => X"10000015",
		16#3db7# => X"a86e0000",
		16#3db8# => X"844b0000",
		16#3db9# => X"d4041000",
		16#3dba# => X"9c400000",
		16#3dbb# => X"d40b1010",
		16#3dbc# => X"d40b100c",
		16#3dbd# => X"9c21000c",
		16#3dbe# => X"8521fffc",
		16#3dbf# => X"8441fff4",
		16#3dc0# => X"44004800",
		16#3dc1# => X"85c1fff8",
		16#3dc2# => X"9c800004",
		16#3dc3# => X"04000c14",
		16#3dc4# => X"9ca00021",
		16#3dc5# => X"a88b0000",
		16#3dc6# => X"bc040000",
		16#3dc7# => X"0fffffeb",
		16#3dc8# => X"d40e584c",
		16#3dc9# => X"03fffff5",
		16#3dca# => X"9c21000c",
		16#3dcb# => X"9c800001",
		16#3dcc# => X"e1c41008",
		16#3dcd# => X"9cae0005",
		16#3dce# => X"04000c09",
		16#3dcf# => X"b8a50002",
		16#3dd0# => X"bc0b0000",
		16#3dd1# => X"13ffffec",
		16#3dd2# => X"15000000",
		16#3dd3# => X"d40b1004",
		16#3dd4# => X"03ffffe6",
		16#3dd5# => X"d40b7008",
		16#3dd6# => X"bc040000",
		16#3dd7# => X"10000009",
		16#3dd8# => X"15000000",
		16#3dd9# => X"84c40004",
		16#3dda# => X"84a3004c",
		16#3ddb# => X"b8660002",
		16#3ddc# => X"e0651800",
		16#3ddd# => X"84a30000",
		16#3dde# => X"d4042800",
		16#3ddf# => X"d4032000",
		16#3de0# => X"44004800",
		16#3de1# => X"15000000",
		16#3de2# => X"d7e117e8",
		16#3de3# => X"d7e177ec",
		16#3de4# => X"d7e187f0",
		16#3de5# => X"d7e197f4",
		16#3de6# => X"d7e14ffc",
		16#3de7# => X"d7e1a7f8",
		16#3de8# => X"a9c40000",
		16#3de9# => X"9c21ffe8",
		16#3dea# => X"aa430000",
		16#3deb# => X"a8460000",
		16#3dec# => X"86040010",
		16#3ded# => X"9ce40014",
		16#3dee# => X"9d000000",
		16#3def# => X"84870000",
		16#3df0# => X"9d080001",
		16#3df1# => X"a4c4ffff",
		16#3df2# => X"b8840050",
		16#3df3# => X"e0c53306",
		16#3df4# => X"e0852306",
		16#3df5# => X"e0c23000",
		16#3df6# => X"e5504000",
		16#3df7# => X"b8460050",
		16#3df8# => X"a4c6ffff",
		16#3df9# => X"e0422000",
		16#3dfa# => X"b8820010",
		16#3dfb# => X"b8420050",
		16#3dfc# => X"e0c43000",
		16#3dfd# => X"d4073000",
		16#3dfe# => X"13fffff1",
		16#3dff# => X"9ce70004",
		16#3e00# => X"bc020000",
		16#3e01# => X"1000000c",
		16#3e02# => X"15000000",
		16#3e03# => X"846e0008",
		16#3e04# => X"e5901800",
		16#3e05# => X"0c000011",
		16#3e06# => X"a8720000",
		16#3e07# => X"9c700005",
		16#3e08# => X"9e100001",
		16#3e09# => X"b8630002",
		16#3e0a# => X"d40e8010",
		16#3e0b# => X"e06e1800",
		16#3e0c# => X"d4031000",
		16#3e0d# => X"9c210018",
		16#3e0e# => X"a96e0000",
		16#3e0f# => X"8521fffc",
		16#3e10# => X"8441ffe8",
		16#3e11# => X"85c1ffec",
		16#3e12# => X"8601fff0",
		16#3e13# => X"8641fff4",
		16#3e14# => X"44004800",
		16#3e15# => X"8681fff8",
		16#3e16# => X"848e0004",
		16#3e17# => X"07ffff92",
		16#3e18# => X"9c840001",
		16#3e19# => X"84ae0010",
		16#3e1a# => X"9c8e000c",
		16#3e1b# => X"9ca50002",
		16#3e1c# => X"9c6b000c",
		16#3e1d# => X"b8a50002",
		16#3e1e# => X"07fffe98",
		16#3e1f# => X"aa8b0000",
		16#3e20# => X"846e0004",
		16#3e21# => X"8492004c",
		16#3e22# => X"b8630002",
		16#3e23# => X"e0641800",
		16#3e24# => X"84830000",
		16#3e25# => X"d40e2000",
		16#3e26# => X"d4037000",
		16#3e27# => X"03ffffe0",
		16#3e28# => X"a9d40000",
		16#3e29# => X"d7e177e8",
		16#3e2a# => X"d7e187ec",
		16#3e2b# => X"d7e197f0",
		16#3e2c# => X"d7e1a7f4",
		16#3e2d# => X"d7e1b7f8",
		16#3e2e# => X"d7e14ffc",
		16#3e2f# => X"d7e117e4",
		16#3e30# => X"a9c30000",
		16#3e31# => X"9c21ffe4",
		16#3e32# => X"aa840000",
		16#3e33# => X"9c660008",
		16#3e34# => X"9c800009",
		16#3e35# => X"aa060000",
		16#3e36# => X"aa450000",
		16#3e37# => X"07ffd4c9",
		16#3e38# => X"aac70000",
		16#3e39# => X"bdab0001",
		16#3e3a# => X"10000007",
		16#3e3b# => X"9c800000",
		16#3e3c# => X"9c400001",
		16#3e3d# => X"e0421000",
		16#3e3e# => X"e54b1000",
		16#3e3f# => X"13fffffe",
		16#3e40# => X"9c840001",
		16#3e41# => X"a86e0000",
		16#3e42# => X"07ffff67",
		16#3e43# => X"9c400001",
		16#3e44# => X"d40bb014",
		16#3e45# => X"bdb20009",
		16#3e46# => X"10000029",
		16#3e47# => X"d40b1010",
		16#3e48# => X"9ed40009",
		16#3e49# => X"9c400009",
		16#3e4a# => X"e0941000",
		16#3e4b# => X"a86e0000",
		16#3e4c# => X"90c40000",
		16#3e4d# => X"9ca0000a",
		16#3e4e# => X"a88b0000",
		16#3e4f# => X"9cc6ffd0",
		16#3e50# => X"07ffff92",
		16#3e51# => X"9c420001",
		16#3e52# => X"e5521000",
		16#3e53# => X"13fffff8",
		16#3e54# => X"e0941000",
		16#3e55# => X"e2969000",
		16#3e56# => X"9e94fff8",
		16#3e57# => X"e5b09000",
		16#3e58# => X"1000000e",
		16#3e59# => X"9c400000",
		16#3e5a# => X"e0941000",
		16#3e5b# => X"a86e0000",
		16#3e5c# => X"90e40000",
		16#3e5d# => X"9ca0000a",
		16#3e5e# => X"a88b0000",
		16#3e5f# => X"9cc7ffd0",
		16#3e60# => X"07ffff82",
		16#3e61# => X"9c420001",
		16#3e62# => X"e0629000",
		16#3e63# => X"e5501800",
		16#3e64# => X"13fffff7",
		16#3e65# => X"e0941000",
		16#3e66# => X"9c21001c",
		16#3e67# => X"8521fffc",
		16#3e68# => X"8441ffe4",
		16#3e69# => X"85c1ffe8",
		16#3e6a# => X"8601ffec",
		16#3e6b# => X"8641fff0",
		16#3e6c# => X"8681fff4",
		16#3e6d# => X"44004800",
		16#3e6e# => X"86c1fff8",
		16#3e6f# => X"9e94000a",
		16#3e70# => X"03ffffe7",
		16#3e71# => X"9e400009",
		16#3e72# => X"d7e117fc",
		16#3e73# => X"1840ffff",
		16#3e74# => X"9d600000",
		16#3e75# => X"e0831003",
		16#3e76# => X"e4245800",
		16#3e77# => X"10000004",
		16#3e78# => X"9c21fffc",
		16#3e79# => X"b8630010",
		16#3e7a# => X"9d600010",
		16#3e7b# => X"1840ff00",
		16#3e7c# => X"e0831003",
		16#3e7d# => X"bc240000",
		16#3e7e# => X"10000004",
		16#3e7f# => X"1840f000",
		16#3e80# => X"b8630008",
		16#3e81# => X"9d6b0008",
		16#3e82# => X"e0831003",
		16#3e83# => X"bc240000",
		16#3e84# => X"10000004",
		16#3e85# => X"1840c000",
		16#3e86# => X"b8630004",
		16#3e87# => X"9d6b0004",
		16#3e88# => X"e0831003",
		16#3e89# => X"bc240000",
		16#3e8a# => X"10000005",
		16#3e8b# => X"bd830000",
		16#3e8c# => X"b8630002",
		16#3e8d# => X"9d6b0002",
		16#3e8e# => X"bd830000",
		16#3e8f# => X"10000007",
		16#3e90# => X"15000000",
		16#3e91# => X"18404000",
		16#3e92# => X"e0631003",
		16#3e93# => X"bc030000",
		16#3e94# => X"10000005",
		16#3e95# => X"9d6b0001",
		16#3e96# => X"9c210004",
		16#3e97# => X"44004800",
		16#3e98# => X"8441fffc",
		16#3e99# => X"9c210004",
		16#3e9a# => X"9d600020",
		16#3e9b# => X"44004800",
		16#3e9c# => X"8441fffc",
		16#3e9d# => X"84830000",
		16#3e9e# => X"a5640007",
		16#3e9f# => X"bc0b0000",
		16#3ea0# => X"1000000e",
		16#3ea1# => X"a4a4ffff",
		16#3ea2# => X"a4a40001",
		16#3ea3# => X"9d600000",
		16#3ea4# => X"e4255800",
		16#3ea5# => X"10000007",
		16#3ea6# => X"a4a40002",
		16#3ea7# => X"e4055800",
		16#3ea8# => X"0c00002a",
		16#3ea9# => X"9d600002",
		16#3eaa# => X"b8840042",
		16#3eab# => X"d4032000",
		16#3eac# => X"44004800",
		16#3ead# => X"15000000",
		16#3eae# => X"bc250000",
		16#3eaf# => X"10000005",
		16#3eb0# => X"a4a400ff",
		16#3eb1# => X"b8840050",
		16#3eb2# => X"9d600010",
		16#3eb3# => X"a4a400ff",
		16#3eb4# => X"bc250000",
		16#3eb5# => X"10000005",
		16#3eb6# => X"a4a4000f",
		16#3eb7# => X"b8840048",
		16#3eb8# => X"9d6b0008",
		16#3eb9# => X"a4a4000f",
		16#3eba# => X"bc250000",
		16#3ebb# => X"10000005",
		16#3ebc# => X"a4a40003",
		16#3ebd# => X"b8840044",
		16#3ebe# => X"9d6b0004",
		16#3ebf# => X"a4a40003",
		16#3ec0# => X"bc250000",
		16#3ec1# => X"10000005",
		16#3ec2# => X"a4a40001",
		16#3ec3# => X"b8840042",
		16#3ec4# => X"9d6b0002",
		16#3ec5# => X"a4a40001",
		16#3ec6# => X"bc250000",
		16#3ec7# => X"10000007",
		16#3ec8# => X"15000000",
		16#3ec9# => X"b8840041",
		16#3eca# => X"bc040000",
		16#3ecb# => X"10000005",
		16#3ecc# => X"15000000",
		16#3ecd# => X"9d6b0001",
		16#3ece# => X"44004800",
		16#3ecf# => X"d4032000",
		16#3ed0# => X"44004800",
		16#3ed1# => X"9d600020",
		16#3ed2# => X"b8840041",
		16#3ed3# => X"9d600001",
		16#3ed4# => X"44004800",
		16#3ed5# => X"d4032000",
		16#3ed6# => X"d7e14ffc",
		16#3ed7# => X"d7e117f8",
		16#3ed8# => X"a8440000",
		16#3ed9# => X"9c21fff8",
		16#3eda# => X"07fffecf",
		16#3edb# => X"9c800001",
		16#3edc# => X"9c800001",
		16#3edd# => X"d40b1014",
		16#3ede# => X"d40b2010",
		16#3edf# => X"9c210008",
		16#3ee0# => X"8521fffc",
		16#3ee1# => X"44004800",
		16#3ee2# => X"8441fff8",
		16#3ee3# => X"d7e177ec",
		16#3ee4# => X"d7e187f0",
		16#3ee5# => X"d7e197f4",
		16#3ee6# => X"d7e1a7f8",
		16#3ee7# => X"d7e14ffc",
		16#3ee8# => X"d7e117e8",
		16#3ee9# => X"86440010",
		16#3eea# => X"86850010",
		16#3eeb# => X"9c21ffe8",
		16#3eec# => X"a9c40000",
		16#3eed# => X"e572a000",
		16#3eee# => X"10000008",
		16#3eef# => X"aa050000",
		16#3ef0# => X"a8920000",
		16#3ef1# => X"a84e0000",
		16#3ef2# => X"aa540000",
		16#3ef3# => X"a9c50000",
		16#3ef4# => X"aa840000",
		16#3ef5# => X"aa020000",
		16#3ef6# => X"e0549000",
		16#3ef7# => X"84ae0008",
		16#3ef8# => X"e5a22800",
		16#3ef9# => X"10000003",
		16#3efa# => X"848e0004",
		16#3efb# => X"9c840001",
		16#3efc# => X"07fffead",
		16#3efd# => X"15000000",
		16#3efe# => X"9ea20005",
		16#3eff# => X"9e6b0014",
		16#3f00# => X"bab50002",
		16#3f01# => X"e2aba800",
		16#3f02# => X"e473a800",
		16#3f03# => X"10000009",
		16#3f04# => X"9ef40005",
		16#3f05# => X"a8d30000",
		16#3f06# => X"9c600000",
		16#3f07# => X"d4061800",
		16#3f08# => X"9cc60004",
		16#3f09# => X"e4553000",
		16#3f0a# => X"13fffffd",
		16#3f0b# => X"9ef40005",
		16#3f0c# => X"9d920005",
		16#3f0d# => X"baf70002",
		16#3f0e# => X"b98c0002",
		16#3f0f# => X"9e300014",
		16#3f10# => X"e2f0b800",
		16#3f11# => X"9f2e0014",
		16#3f12# => X"e471b800",
		16#3f13# => X"10000045",
		16#3f14# => X"e18e6000",
		16#3f15# => X"84f10000",
		16#3f16# => X"a4a7ffff",
		16#3f17# => X"bc050000",
		16#3f18# => X"1000001e",
		16#3f19# => X"b8e70050",
		16#3f1a# => X"a8730000",
		16#3f1b# => X"a8990000",
		16#3f1c# => X"9cc00000",
		16#3f1d# => X"85a40000",
		16#3f1e# => X"85030000",
		16#3f1f# => X"a4edffff",
		16#3f20# => X"b9ad0050",
		16#3f21# => X"e0e72b06",
		16#3f22# => X"e1ad2b06",
		16#3f23# => X"a5e8ffff",
		16#3f24# => X"b9080050",
		16#3f25# => X"e0e77800",
		16#3f26# => X"9c840004",
		16#3f27# => X"e0e73000",
		16#3f28# => X"e0cd4000",
		16#3f29# => X"b9070050",
		16#3f2a# => X"a4e7ffff",
		16#3f2b# => X"e44c2000",
		16#3f2c# => X"e0c64000",
		16#3f2d# => X"b9060010",
		16#3f2e# => X"b8c60050",
		16#3f2f# => X"e0e83804",
		16#3f30# => X"d4033800",
		16#3f31# => X"13ffffec",
		16#3f32# => X"9c630004",
		16#3f33# => X"d4033000",
		16#3f34# => X"84f10000",
		16#3f35# => X"b8e70050",
		16#3f36# => X"bc070000",
		16#3f37# => X"1000001d",
		16#3f38# => X"a8930000",
		16#3f39# => X"84b30000",
		16#3f3a# => X"a8c50000",
		16#3f3b# => X"a8790000",
		16#3f3c# => X"9d000000",
		16#3f3d# => X"85a30000",
		16#3f3e# => X"b8c60050",
		16#3f3f# => X"a5adffff",
		16#3f40# => X"a4a5ffff",
		16#3f41# => X"e1a76b06",
		16#3f42# => X"e1086800",
		16#3f43# => X"e0c83000",
		16#3f44# => X"b9a60010",
		16#3f45# => X"b9060050",
		16#3f46# => X"e0ad2804",
		16#3f47# => X"d4042800",
		16#3f48# => X"9c840004",
		16#3f49# => X"94a30000",
		16#3f4a# => X"e0a72b06",
		16#3f4b# => X"84c40000",
		16#3f4c# => X"9c630004",
		16#3f4d# => X"a5a6ffff",
		16#3f4e# => X"e44c1800",
		16#3f4f# => X"e0a56800",
		16#3f50# => X"e0a54000",
		16#3f51# => X"13ffffec",
		16#3f52# => X"b9050050",
		16#3f53# => X"d4042800",
		16#3f54# => X"9e310004",
		16#3f55# => X"e4b78800",
		16#3f56# => X"0fffffbf",
		16#3f57# => X"9e730004",
		16#3f58# => X"bda20000",
		16#3f59# => X"10000012",
		16#3f5a# => X"15000000",
		16#3f5b# => X"9c75fffc",
		16#3f5c# => X"84830000",
		16#3f5d# => X"bc240000",
		16#3f5e# => X"0c00000a",
		16#3f5f# => X"9c42ffff",
		16#3f60# => X"9c420001",
		16#3f61# => X"0000000b",
		16#3f62# => X"d40b1010",
		16#3f63# => X"84830000",
		16#3f64# => X"bc040000",
		16#3f65# => X"0c000006",
		16#3f66# => X"15000000",
		16#3f67# => X"9c42ffff",
		16#3f68# => X"bda20000",
		16#3f69# => X"0ffffffa",
		16#3f6a# => X"9c63fffc",
		16#3f6b# => X"d40b1010",
		16#3f6c# => X"9c210018",
		16#3f6d# => X"8521fffc",
		16#3f6e# => X"8441ffe8",
		16#3f6f# => X"85c1ffec",
		16#3f70# => X"8601fff0",
		16#3f71# => X"8641fff4",
		16#3f72# => X"44004800",
		16#3f73# => X"8681fff8",
		16#3f74# => X"d7e117e8",
		16#3f75# => X"d7e187f0",
		16#3f76# => X"d7e1a7f8",
		16#3f77# => X"d7e14ffc",
		16#3f78# => X"d7e177ec",
		16#3f79# => X"d7e197f4",
		16#3f7a# => X"a8450000",
		16#3f7b# => X"a4a50003",
		16#3f7c# => X"9c21ffe8",
		16#3f7d# => X"aa830000",
		16#3f7e# => X"bc050000",
		16#3f7f# => X"0c00003c",
		16#3f80# => X"aa040000",
		16#3f81# => X"b8420082",
		16#3f82# => X"bc020000",
		16#3f83# => X"10000026",
		16#3f84# => X"15000000",
		16#3f85# => X"85d40048",
		16#3f86# => X"bc2e0000",
		16#3f87# => X"1000000e",
		16#3f88# => X"a4820001",
		16#3f89# => X"0000003c",
		16#3f8a# => X"a8740000",
		16#3f8b# => X"b8420081",
		16#3f8c# => X"bc020000",
		16#3f8d# => X"1000001c",
		16#3f8e# => X"15000000",
		16#3f8f# => X"864e0000",
		16#3f90# => X"bc320000",
		16#3f91# => X"0c000021",
		16#3f92# => X"a88e0000",
		16#3f93# => X"a9d20000",
		16#3f94# => X"a4820001",
		16#3f95# => X"bc040000",
		16#3f96# => X"13fffff5",
		16#3f97# => X"a8900000",
		16#3f98# => X"a8ae0000",
		16#3f99# => X"07ffff4a",
		16#3f9a# => X"a8740000",
		16#3f9b# => X"bc100000",
		16#3f9c# => X"1000001d",
		16#3f9d# => X"15000000",
		16#3f9e# => X"84700004",
		16#3f9f# => X"8494004c",
		16#3fa0# => X"b8630002",
		16#3fa1# => X"b8420081",
		16#3fa2# => X"e0641800",
		16#3fa3# => X"bc020000",
		16#3fa4# => X"84830000",
		16#3fa5# => X"d4102000",
		16#3fa6# => X"d4038000",
		16#3fa7# => X"0fffffe8",
		16#3fa8# => X"aa0b0000",
		16#3fa9# => X"9c210018",
		16#3faa# => X"a9700000",
		16#3fab# => X"8521fffc",
		16#3fac# => X"8441ffe8",
		16#3fad# => X"85c1ffec",
		16#3fae# => X"8601fff0",
		16#3faf# => X"8641fff4",
		16#3fb0# => X"44004800",
		16#3fb1# => X"8681fff8",
		16#3fb2# => X"a8ae0000",
		16#3fb3# => X"07ffff30",
		16#3fb4# => X"a8740000",
		16#3fb5# => X"d40e5800",
		16#3fb6# => X"d40b9000",
		16#3fb7# => X"03ffffdd",
		16#3fb8# => X"a9cb0000",
		16#3fb9# => X"03ffffd2",
		16#3fba# => X"aa0b0000",
		16#3fbb# => X"9ca5ffff",
		16#3fbc# => X"18e00001",
		16#3fbd# => X"b8a50002",
		16#3fbe# => X"a8e74230",
		16#3fbf# => X"9cc00000",
		16#3fc0# => X"e0a53800",
		16#3fc1# => X"07fffe21",
		16#3fc2# => X"84a50000",
		16#3fc3# => X"03ffffbe",
		16#3fc4# => X"aa0b0000",
		16#3fc5# => X"07ffff11",
		16#3fc6# => X"9c800271",
		16#3fc7# => X"9c600000",
		16#3fc8# => X"d4145848",
		16#3fc9# => X"a9cb0000",
		16#3fca# => X"03ffffca",
		16#3fcb# => X"d40b1800",
		16#3fcc# => X"d7e177ec",
		16#3fcd# => X"85c40010",
		16#3fce# => X"d7e187f0",
		16#3fcf# => X"ba050085",
		16#3fd0# => X"9dce0001",
		16#3fd1# => X"d7e117e8",
		16#3fd2# => X"d7e197f4",
		16#3fd3# => X"d7e1a7f8",
		16#3fd4# => X"84c40008",
		16#3fd5# => X"d7e14ffc",
		16#3fd6# => X"e1ce8000",
		16#3fd7# => X"a8440000",
		16#3fd8# => X"9c21ffe8",
		16#3fd9# => X"aa850000",
		16#3fda# => X"aa430000",
		16#3fdb# => X"e5ae3000",
		16#3fdc# => X"10000006",
		16#3fdd# => X"84840004",
		16#3fde# => X"e0c63000",
		16#3fdf# => X"e54e3000",
		16#3fe0# => X"13fffffe",
		16#3fe1# => X"9c840001",
		16#3fe2# => X"07fffdc7",
		16#3fe3# => X"a8720000",
		16#3fe4# => X"bdb00000",
		16#3fe5# => X"a90b0000",
		16#3fe6# => X"1000000c",
		16#3fe7# => X"9ccb0014",
		16#3fe8# => X"9ce00000",
		16#3fe9# => X"9c600000",
		16#3fea# => X"9ce70001",
		16#3feb# => X"d4061800",
		16#3fec# => X"e4278000",
		16#3fed# => X"13fffffd",
		16#3fee# => X"9cc60004",
		16#3fef# => X"9cc70005",
		16#3ff0# => X"b8c60002",
		16#3ff1# => X"e0c83000",
		16#3ff2# => X"85620010",
		16#3ff3# => X"a4b4001f",
		16#3ff4# => X"9d6b0005",
		16#3ff5# => X"9ce20014",
		16#3ff6# => X"b96b0002",
		16#3ff7# => X"bc050000",
		16#3ff8# => X"10000025",
		16#3ff9# => X"e1625800",
		16#3ffa# => X"9da00020",
		16#3ffb# => X"9c800000",
		16#3ffc# => X"e1ad2802",
		16#3ffd# => X"85870000",
		16#3ffe# => X"e18c2808",
		16#3fff# => X"e0846004",
		16#4000# => X"d4062000",
		16#4001# => X"9cc60004",
		16#4002# => X"84870000",
		16#4003# => X"9ce70004",
		16#4004# => X"e44b3800",
		16#4005# => X"13fffff8",
		16#4006# => X"e0846848",
		16#4007# => X"bc040000",
		16#4008# => X"10000003",
		16#4009# => X"d4062000",
		16#400a# => X"9dce0001",
		16#400b# => X"84620004",
		16#400c# => X"8492004c",
		16#400d# => X"b8630002",
		16#400e# => X"9dceffff",
		16#400f# => X"a9680000",
		16#4010# => X"e0641800",
		16#4011# => X"d4087010",
		16#4012# => X"84830000",
		16#4013# => X"d4022000",
		16#4014# => X"d4031000",
		16#4015# => X"9c210018",
		16#4016# => X"8521fffc",
		16#4017# => X"8441ffe8",
		16#4018# => X"85c1ffec",
		16#4019# => X"8601fff0",
		16#401a# => X"8641fff4",
		16#401b# => X"44004800",
		16#401c# => X"8681fff8",
		16#401d# => X"84670000",
		16#401e# => X"9ce70004",
		16#401f# => X"d4061800",
		16#4020# => X"e44b3800",
		16#4021# => X"0fffffea",
		16#4022# => X"9cc60004",
		16#4023# => X"84670000",
		16#4024# => X"9ce70004",
		16#4025# => X"d4061800",
		16#4026# => X"e44b3800",
		16#4027# => X"13fffff6",
		16#4028# => X"9cc60004",
		16#4029# => X"03ffffe3",
		16#402a# => X"84620004",
		16#402b# => X"85630010",
		16#402c# => X"84a40010",
		16#402d# => X"e16b2802",
		16#402e# => X"bc2b0000",
		16#402f# => X"10000010",
		16#4030# => X"15000000",
		16#4031# => X"9ca50005",
		16#4032# => X"9ce30014",
		16#4033# => X"b8a50002",
		16#4034# => X"e0632800",
		16#4035# => X"e0842800",
		16#4036# => X"9c63fffc",
		16#4037# => X"9c84fffc",
		16#4038# => X"84c30000",
		16#4039# => X"84a40000",
		16#403a# => X"e4062800",
		16#403b# => X"0c000006",
		16#403c# => X"e4871800",
		16#403d# => X"13fffff9",
		16#403e# => X"15000000",
		16#403f# => X"44004800",
		16#4040# => X"15000000",
		16#4041# => X"e4662800",
		16#4042# => X"13fffffd",
		16#4043# => X"9d600001",
		16#4044# => X"44004800",
		16#4045# => X"9d60ffff",
		16#4046# => X"d7e117ec",
		16#4047# => X"a8440000",
		16#4048# => X"d7e177f0",
		16#4049# => X"d7e187f4",
		16#404a# => X"d7e197f8",
		16#404b# => X"d7e14ffc",
		16#404c# => X"aa430000",
		16#404d# => X"9c21ffec",
		16#404e# => X"a8850000",
		16#404f# => X"a8620000",
		16#4050# => X"07ffffdb",
		16#4051# => X"a9c50000",
		16#4052# => X"bc2b0000",
		16#4053# => X"0c00005a",
		16#4054# => X"aa0b0000",
		16#4055# => X"bd8b0000",
		16#4056# => X"10000053",
		16#4057# => X"9e000001",
		16#4058# => X"9e000000",
		16#4059# => X"a8720000",
		16#405a# => X"07fffd4f",
		16#405b# => X"84820004",
		16#405c# => X"846e0010",
		16#405d# => X"85820010",
		16#405e# => X"9c630005",
		16#405f# => X"9dec0005",
		16#4060# => X"b8630002",
		16#4061# => X"b9ef0002",
		16#4062# => X"9cee0014",
		16#4063# => X"d40b800c",
		16#4064# => X"e1ce1800",
		16#4065# => X"9cc20014",
		16#4066# => X"e1e27800",
		16#4067# => X"9c6b0014",
		16#4068# => X"9d000000",
		16#4069# => X"86a60000",
		16#406a# => X"86670000",
		16#406b# => X"a635ffff",
		16#406c# => X"a5b3ffff",
		16#406d# => X"bab50050",
		16#406e# => X"e1b16802",
		16#406f# => X"ba730050",
		16#4070# => X"e1ad4000",
		16#4071# => X"9ce70004",
		16#4072# => X"ba2d0090",
		16#4073# => X"e1159802",
		16#4074# => X"a5adffff",
		16#4075# => X"e1088800",
		16#4076# => X"9cc60004",
		16#4077# => X"ba280010",
		16#4078# => X"e44e3800",
		16#4079# => X"b9080090",
		16#407a# => X"e1b16804",
		16#407b# => X"d4036800",
		16#407c# => X"13ffffed",
		16#407d# => X"9c630004",
		16#407e# => X"a8430000",
		16#407f# => X"e4af3000",
		16#4080# => X"10000017",
		16#4081# => X"a8860000",
		16#4082# => X"84e60000",
		16#4083# => X"9cc60004",
		16#4084# => X"a4a7ffff",
		16#4085# => X"b8e70050",
		16#4086# => X"e0a82800",
		16#4087# => X"e44f3000",
		16#4088# => X"b9050090",
		16#4089# => X"a4a5ffff",
		16#408a# => X"e1083800",
		16#408b# => X"b8e80010",
		16#408c# => X"b9080090",
		16#408d# => X"e0a72804",
		16#408e# => X"d4032800",
		16#408f# => X"13fffff3",
		16#4090# => X"9c630004",
		16#4091# => X"ac64ffff",
		16#4092# => X"9c80fffc",
		16#4093# => X"e0637800",
		16#4094# => X"e0632003",
		16#4095# => X"9c630004",
		16#4096# => X"e0621800",
		16#4097# => X"9c63fffc",
		16#4098# => X"84430000",
		16#4099# => X"bc220000",
		16#409a# => X"10000007",
		16#409b# => X"15000000",
		16#409c# => X"9c63fffc",
		16#409d# => X"84430000",
		16#409e# => X"bc020000",
		16#409f# => X"13fffffd",
		16#40a0# => X"9d8cffff",
		16#40a1# => X"d40b6010",
		16#40a2# => X"9c210014",
		16#40a3# => X"8521fffc",
		16#40a4# => X"8441ffec",
		16#40a5# => X"85c1fff0",
		16#40a6# => X"8601fff4",
		16#40a7# => X"44004800",
		16#40a8# => X"8641fff8",
		16#40a9# => X"a8620000",
		16#40aa# => X"a84e0000",
		16#40ab# => X"03ffffae",
		16#40ac# => X"a9c30000",
		16#40ad# => X"a8720000",
		16#40ae# => X"9c400001",
		16#40af# => X"07fffcfa",
		16#40b0# => X"a88b0000",
		16#40b1# => X"d40b8014",
		16#40b2# => X"d40b1010",
		16#40b3# => X"9c210014",
		16#40b4# => X"8521fffc",
		16#40b5# => X"8441ffec",
		16#40b6# => X"85c1fff0",
		16#40b7# => X"8601fff4",
		16#40b8# => X"44004800",
		16#40b9# => X"8641fff8",
		16#40ba# => X"d7e117fc",
		16#40bb# => X"18407ff0",
		16#40bc# => X"9c21fffc",
		16#40bd# => X"e0631003",
		16#40be# => X"1840fcc0",
		16#40bf# => X"e0631000",
		16#40c0# => X"bda30000",
		16#40c1# => X"10000007",
		16#40c2# => X"9c800000",
		16#40c3# => X"9c210004",
		16#40c4# => X"a9630000",
		16#40c5# => X"a9840000",
		16#40c6# => X"44004800",
		16#40c7# => X"8441fffc",
		16#40c8# => X"e0601802",
		16#40c9# => X"b8630094",
		16#40ca# => X"bd430013",
		16#40cb# => X"0c00000e",
		16#40cc# => X"9ca3ffec",
		16#40cd# => X"9c800001",
		16#40ce# => X"bd45001e",
		16#40cf# => X"13fffff4",
		16#40d0# => X"9c600000",
		16#40d1# => X"9cc0001f",
		16#40d2# => X"9c210004",
		16#40d3# => X"e0a62802",
		16#40d4# => X"a9630000",
		16#40d5# => X"e0842808",
		16#40d6# => X"8441fffc",
		16#40d7# => X"44004800",
		16#40d8# => X"a9840000",
		16#40d9# => X"18a00008",
		16#40da# => X"9c800000",
		16#40db# => X"e0651888",
		16#40dc# => X"9c210004",
		16#40dd# => X"a9840000",
		16#40de# => X"a9630000",
		16#40df# => X"44004800",
		16#40e0# => X"8441fffc",
		16#40e1# => X"d7e197f4",
		16#40e2# => X"86430010",
		16#40e3# => X"d7e117e8",
		16#40e4# => X"9e520005",
		16#40e5# => X"d7e177ec",
		16#40e6# => X"ba520002",
		16#40e7# => X"d7e187f0",
		16#40e8# => X"d7e1a7f8",
		16#40e9# => X"e2439000",
		16#40ea# => X"d7e14ffc",
		16#40eb# => X"9c52fffc",
		16#40ec# => X"9c21ffe8",
		16#40ed# => X"85c20000",
		16#40ee# => X"9e030014",
		16#40ef# => X"a86e0000",
		16#40f0# => X"07fffd82",
		16#40f1# => X"aa840000",
		16#40f2# => X"9c600020",
		16#40f3# => X"bd4b000a",
		16#40f4# => X"e0635802",
		16#40f5# => X"10000019",
		16#40f6# => X"d4141800",
		16#40f7# => X"9ca0000b",
		16#40f8# => X"18c03ff0",
		16#40f9# => X"e0a55802",
		16#40fa# => X"9c800000",
		16#40fb# => X"e06e2848",
		16#40fc# => X"e4701000",
		16#40fd# => X"10000004",
		16#40fe# => X"e0633004",
		16#40ff# => X"8482fffc",
		16#4100# => X"e0842848",
		16#4101# => X"9d6b0015",
		16#4102# => X"e1ce5808",
		16#4103# => X"e1c47004",
		16#4104# => X"9c210018",
		16#4105# => X"a98e0000",
		16#4106# => X"8521fffc",
		16#4107# => X"a9630000",
		16#4108# => X"8441ffe8",
		16#4109# => X"85c1ffec",
		16#410a# => X"8601fff0",
		16#410b# => X"8641fff4",
		16#410c# => X"44004800",
		16#410d# => X"8681fff8",
		16#410e# => X"e4701000",
		16#410f# => X"10000004",
		16#4110# => X"9c800000",
		16#4111# => X"9c52fff8",
		16#4112# => X"84820000",
		16#4113# => X"9d6bfff5",
		16#4114# => X"bc0b0000",
		16#4115# => X"10000010",
		16#4116# => X"19003ff0",
		16#4117# => X"9cc00020",
		16#4118# => X"e06e5808",
		16#4119# => X"e0c65802",
		16#411a# => X"e0e43048",
		16#411b# => X"e0634004",
		16#411c# => X"9ca00000",
		16#411d# => X"e4a28000",
		16#411e# => X"10000004",
		16#411f# => X"e0633804",
		16#4120# => X"84a2fffc",
		16#4121# => X"e0a53048",
		16#4122# => X"e1c45808",
		16#4123# => X"03ffffe1",
		16#4124# => X"e1c57004",
		16#4125# => X"18403ff0",
		16#4126# => X"e06e1004",
		16#4127# => X"03ffffdd",
		16#4128# => X"a9c40000",
		16#4129# => X"d7e117e4",
		16#412a# => X"d7e177e8",
		16#412b# => X"d7e187ec",
		16#412c# => X"d7e197f0",
		16#412d# => X"d7e1a7f4",
		16#412e# => X"d7e1b7f8",
		16#412f# => X"aa040000",
		16#4130# => X"d7e14ffc",
		16#4131# => X"9c800001",
		16#4132# => X"9c21ffdc",
		16#4133# => X"aac60000",
		16#4134# => X"aa870000",
		16#4135# => X"07fffc74",
		16#4136# => X"aa450000",
		16#4137# => X"18607fff",
		16#4138# => X"a84b0000",
		16#4139# => X"a863ffff",
		16#413a# => X"e1d01803",
		16#413b# => X"1860000f",
		16#413c# => X"b9ce0054",
		16#413d# => X"a863ffff",
		16#413e# => X"e2101803",
		16#413f# => X"bc0e0000",
		16#4140# => X"10000005",
		16#4141# => X"d4018000",
		16#4142# => X"18600010",
		16#4143# => X"e2101804",
		16#4144# => X"d4018000",
		16#4145# => X"bc120000",
		16#4146# => X"1000001a",
		16#4147# => X"a8610000",
		16#4148# => X"9c610004",
		16#4149# => X"07fffd54",
		16#414a# => X"d4019004",
		16#414b# => X"bc0b0000",
		16#414c# => X"0c000030",
		16#414d# => X"9c800020",
		16#414e# => X"84810004",
		16#414f# => X"84610000",
		16#4150# => X"d4022014",
		16#4151# => X"d4021818",
		16#4152# => X"bc030000",
		16#4153# => X"10000003",
		16#4154# => X"9e000001",
		16#4155# => X"9e000002",
		16#4156# => X"bc0e0000",
		16#4157# => X"10000011",
		16#4158# => X"d4028010",
		16#4159# => X"9dcefbcd",
		16#415a# => X"9c600035",
		16#415b# => X"e1ce5800",
		16#415c# => X"e1635802",
		16#415d# => X"d4167000",
		16#415e# => X"00000014",
		16#415f# => X"d4145800",
		16#4160# => X"07fffd3d",
		16#4161# => X"9e000001",
		16#4162# => X"84610000",
		16#4163# => X"d4028010",
		16#4164# => X"d4021814",
		16#4165# => X"bc0e0000",
		16#4166# => X"0ffffff3",
		16#4167# => X"9d6b0020",
		16#4168# => X"9c700004",
		16#4169# => X"9d6bfbce",
		16#416a# => X"b8630002",
		16#416b# => X"ba100005",
		16#416c# => X"d4165800",
		16#416d# => X"e0621800",
		16#416e# => X"07fffd04",
		16#416f# => X"84630000",
		16#4170# => X"e1705802",
		16#4171# => X"d4145800",
		16#4172# => X"9c210024",
		16#4173# => X"a9620000",
		16#4174# => X"8521fffc",
		16#4175# => X"8441ffe4",
		16#4176# => X"85c1ffe8",
		16#4177# => X"8601ffec",
		16#4178# => X"8641fff0",
		16#4179# => X"8681fff4",
		16#417a# => X"44004800",
		16#417b# => X"86c1fff8",
		16#417c# => X"84610000",
		16#417d# => X"e0845802",
		16#417e# => X"84a10004",
		16#417f# => X"e0832008",
		16#4180# => X"e0635848",
		16#4181# => X"e0842804",
		16#4182# => X"d4011800",
		16#4183# => X"03ffffce",
		16#4184# => X"d4022014",
		16#4185# => X"d7e14ffc",
		16#4186# => X"d7e117e4",
		16#4187# => X"d7e177e8",
		16#4188# => X"d7e187ec",
		16#4189# => X"d7e197f0",
		16#418a# => X"d7e1a7f4",
		16#418b# => X"d7e1b7f8",
		16#418c# => X"9c21ffdc",
		16#418d# => X"aa440000",
		16#418e# => X"9c810004",
		16#418f# => X"07ffff52",
		16#4190# => X"aa830000",
		16#4191# => X"a8720000",
		16#4192# => X"a8810000",
		16#4193# => X"a9cb0000",
		16#4194# => X"07ffff4d",
		16#4195# => X"aa0c0000",
		16#4196# => X"84740010",
		16#4197# => X"84920010",
		16#4198# => X"84a10004",
		16#4199# => X"e0832002",
		16#419a# => X"84610000",
		16#419b# => X"b8840005",
		16#419c# => X"e0651802",
		16#419d# => X"a84b0000",
		16#419e# => X"e0632000",
		16#419f# => X"aace0000",
		16#41a0# => X"a8ec0000",
		16#41a1# => X"bda30000",
		16#41a2# => X"10000016",
		16#41a3# => X"a8a20000",
		16#41a4# => X"b9c30014",
		16#41a5# => X"e1ceb000",
		16#41a6# => X"a86e0000",
		16#41a7# => X"a8a20000",
		16#41a8# => X"a8900000",
		16#41a9# => X"07ffd933",
		16#41aa# => X"a8c70000",
		16#41ab# => X"9c210024",
		16#41ac# => X"a84b0000",
		16#41ad# => X"a86c0000",
		16#41ae# => X"8521fffc",
		16#41af# => X"e1620004",
		16#41b0# => X"e1830004",
		16#41b1# => X"85c1ffe8",
		16#41b2# => X"8441ffe4",
		16#41b3# => X"8601ffec",
		16#41b4# => X"8641fff0",
		16#41b5# => X"8681fff4",
		16#41b6# => X"44004800",
		16#41b7# => X"86c1fff8",
		16#41b8# => X"b8430014",
		16#41b9# => X"03ffffed",
		16#41ba# => X"e0451002",
		16#41bb# => X"d7e117f8",
		16#41bc# => X"d7e14ffc",
		16#41bd# => X"a8430000",
		16#41be# => X"bd430017",
		16#41bf# => X"0c000017",
		16#41c0# => X"9c21fff8",
		16#41c1# => X"19603ff0",
		16#41c2# => X"9d800000",
		16#41c3# => X"18e00001",
		16#41c4# => X"a86b0000",
		16#41c5# => X"a8e74110",
		16#41c6# => X"a88c0000",
		16#41c7# => X"84a70000",
		16#41c8# => X"84c70004",
		16#41c9# => X"07ffd810",
		16#41ca# => X"9c42ffff",
		16#41cb# => X"bc220000",
		16#41cc# => X"13fffff8",
		16#41cd# => X"18e00001",
		16#41ce# => X"9c210008",
		16#41cf# => X"a84b0000",
		16#41d0# => X"a86c0000",
		16#41d1# => X"8521fffc",
		16#41d2# => X"e1620004",
		16#41d3# => X"e1830004",
		16#41d4# => X"44004800",
		16#41d5# => X"8441fff8",
		16#41d6# => X"b8430003",
		16#41d7# => X"18600001",
		16#41d8# => X"9c210008",
		16#41d9# => X"a8634118",
		16#41da# => X"8521fffc",
		16#41db# => X"e0421800",
		16#41dc# => X"85820004",
		16#41dd# => X"85620000",
		16#41de# => X"a86c0000",
		16#41df# => X"a84b0000",
		16#41e0# => X"e1620004",
		16#41e1# => X"e1830004",
		16#41e2# => X"44004800",
		16#41e3# => X"8441fff8",
		16#41e4# => X"9c84ffff",
		16#41e5# => X"84e50010",
		16#41e6# => X"b9040085",
		16#41e7# => X"9ce70005",
		16#41e8# => X"d7e117fc",
		16#41e9# => X"9d080001",
		16#41ea# => X"b8e70002",
		16#41eb# => X"b9080002",
		16#41ec# => X"9c850014",
		16#41ed# => X"e0e53800",
		16#41ee# => X"9c21fffc",
		16#41ef# => X"e4643800",
		16#41f0# => X"1000000f",
		16#41f1# => X"e1034000",
		16#41f2# => X"a8c30000",
		16#41f3# => X"85640000",
		16#41f4# => X"9c840004",
		16#41f5# => X"d4065800",
		16#41f6# => X"e4472000",
		16#41f7# => X"13fffffc",
		16#41f8# => X"9cc60004",
		16#41f9# => X"e0872802",
		16#41fa# => X"9c40fffc",
		16#41fb# => X"9c84ffeb",
		16#41fc# => X"e0841003",
		16#41fd# => X"9c840004",
		16#41fe# => X"e0632000",
		16#41ff# => X"e4a81800",
		16#4200# => X"10000008",
		16#4201# => X"15000000",
		16#4202# => X"9c400000",
		16#4203# => X"d4031000",
		16#4204# => X"9c630004",
		16#4205# => X"e4481800",
		16#4206# => X"13fffffd",
		16#4207# => X"15000000",
		16#4208# => X"9c210004",
		16#4209# => X"44004800",
		16#420a# => X"8441fffc",
		16#420b# => X"b8a40085",
		16#420c# => X"84c30010",
		16#420d# => X"e5662800",
		16#420e# => X"10000019",
		16#420f# => X"e5462800",
		16#4210# => X"a8a60000",
		16#4211# => X"9ca50005",
		16#4212# => X"9c830014",
		16#4213# => X"b8a50002",
		16#4214# => X"e0632800",
		16#4215# => X"e4641800",
		16#4216# => X"1000000f",
		16#4217# => X"9d600000",
		16#4218# => X"9c63fffc",
		16#4219# => X"84a30000",
		16#421a# => X"bc250000",
		16#421b# => X"1000000a",
		16#421c# => X"9d600001",
		16#421d# => X"e4841800",
		16#421e# => X"0c000018",
		16#421f# => X"9c63fffc",
		16#4220# => X"84a30000",
		16#4221# => X"bc250000",
		16#4222# => X"0ffffffc",
		16#4223# => X"e4841800",
		16#4224# => X"9d600001",
		16#4225# => X"44004800",
		16#4226# => X"15000000",
		16#4227# => X"0fffffea",
		16#4228# => X"a484001f",
		16#4229# => X"bc240000",
		16#422a# => X"0fffffe7",
		16#422b# => X"9cc50005",
		16#422c# => X"b8c60002",
		16#422d# => X"e0c33000",
		16#422e# => X"84c60000",
		16#422f# => X"e0e62048",
		16#4230# => X"e0872008",
		16#4231# => X"e4243000",
		16#4232# => X"0fffffdf",
		16#4233# => X"9d600001",
		16#4234# => X"44004800",
		16#4235# => X"15000000",
		16#4236# => X"44004800",
		16#4237# => X"9d600000",
		16#4238# => X"d7e187dc",
		16#4239# => X"d7e197e0",
		16#423a# => X"d7e1c7ec",
		16#423b# => X"d7e14ffc",
		16#423c# => X"d7e117d4",
		16#423d# => X"d7e177d8",
		16#423e# => X"d7e1a7e4",
		16#423f# => X"d7e1b7e8",
		16#4240# => X"d7e1d7f0",
		16#4241# => X"d7e1e7f4",
		16#4242# => X"d7e1f7f8",
		16#4243# => X"aa040000",
		16#4244# => X"9c21ffd4",
		16#4245# => X"ab030000",
		16#4246# => X"bc240000",
		16#4247# => X"0c00010f",
		16#4248# => X"aa450000",
		16#4249# => X"9c50fff8",
		16#424a# => X"07ffde60",
		16#424b# => X"9dd2000b",
		16#424c# => X"bcae0016",
		16#424d# => X"0c000065",
		16#424e# => X"84c20004",
		16#424f# => X"9c600010",
		16#4250# => X"9c800000",
		16#4251# => X"a9c30000",
		16#4252# => X"e48e9000",
		16#4253# => X"10000003",
		16#4254# => X"9ca00001",
		16#4255# => X"9ca00000",
		16#4256# => X"a4a500ff",
		16#4257# => X"bc250000",
		16#4258# => X"1000010c",
		16#4259# => X"bc040000",
		16#425a# => X"0c00010a",
		16#425b# => X"9ca0fffc",
		16#425c# => X"e2862803",
		16#425d# => X"e5741800",
		16#425e# => X"10000059",
		16#425f# => X"aad40000",
		16#4260# => X"1b800001",
		16#4261# => X"e0e2a000",
		16#4262# => X"ab9c6808",
		16#4263# => X"84bc0008",
		16#4264# => X"e4053800",
		16#4265# => X"10000103",
		16#4266# => X"9d80fffe",
		16#4267# => X"85070004",
		16#4268# => X"e1686003",
		16#4269# => X"e1675800",
		16#426a# => X"856b0004",
		16#426b# => X"a56b0001",
		16#426c# => X"bc0b0000",
		16#426d# => X"10000066",
		16#426e# => X"9d60fffc",
		16#426f# => X"a8e40000",
		16#4270# => X"a4c60001",
		16#4271# => X"bc260000",
		16#4272# => X"1000007a",
		16#4273# => X"9d60fffc",
		16#4274# => X"87420000",
		16#4275# => X"e342d002",
		16#4276# => X"bc070000",
		16#4277# => X"87da0004",
		16#4278# => X"100000ad",
		16#4279# => X"e3de5803",
		16#427a# => X"e4272800",
		16#427b# => X"0c00010f",
		16#427c# => X"9cae0010",
		16#427d# => X"e3dea000",
		16#427e# => X"e2c4f000",
		16#427f# => X"e543b000",
		16#4280# => X"100000a7",
		16#4281# => X"e543f000",
		16#4282# => X"8447000c",
		16#4283# => X"84670008",
		16#4284# => X"9cb4fffc",
		16#4285# => X"d403100c",
		16#4286# => X"d4021808",
		16#4287# => X"845a000c",
		16#4288# => X"847a0008",
		16#4289# => X"9e5a0008",
		16#428a# => X"d403100c",
		16#428b# => X"bc450024",
		16#428c# => X"1000013f",
		16#428d# => X"d4021808",
		16#428e# => X"bca50013",
		16#428f# => X"10000018",
		16#4290# => X"a8520000",
		16#4291# => X"84700000",
		16#4292# => X"9c5a0010",
		16#4293# => X"d4121800",
		16#4294# => X"bca5001b",
		16#4295# => X"84700004",
		16#4296# => X"9e100008",
		16#4297# => X"10000010",
		16#4298# => X"d41a180c",
		16#4299# => X"84700000",
		16#429a# => X"bc250024",
		16#429b# => X"d4021800",
		16#429c# => X"9c5a0018",
		16#429d# => X"84700004",
		16#429e# => X"9e100008",
		16#429f# => X"10000008",
		16#42a0# => X"d41a1814",
		16#42a1# => X"84700000",
		16#42a2# => X"d4021800",
		16#42a3# => X"9c5a0020",
		16#42a4# => X"84700004",
		16#42a5# => X"9e100008",
		16#42a6# => X"d41a181c",
		16#42a7# => X"84700000",
		16#42a8# => X"9e100004",
		16#42a9# => X"d4021800",
		16#42aa# => X"9c620004",
		16#42ab# => X"84500000",
		16#42ac# => X"d4031000",
		16#42ad# => X"a85a0000",
		16#42ae# => X"84900004",
		16#42af# => X"d4032004",
		16#42b0# => X"00000008",
		16#42b1# => X"84da0004",
		16#42b2# => X"9c60fff8",
		16#42b3# => X"e1ce1803",
		16#42b4# => X"a86e0000",
		16#42b5# => X"03ffff9d",
		16#42b6# => X"b88e005f",
		16#42b7# => X"9e420008",
		16#42b8# => X"e0767002",
		16#42b9# => X"bca3000f",
		16#42ba# => X"0c000024",
		16#42bb# => X"e0827000",
		16#42bc# => X"a4c60001",
		16#42bd# => X"e062b000",
		16#42be# => X"e2c6b004",
		16#42bf# => X"d402b004",
		16#42c0# => X"84430004",
		16#42c1# => X"a8420001",
		16#42c2# => X"d4031004",
		16#42c3# => X"07ffdde9",
		16#42c4# => X"a8780000",
		16#42c5# => X"9c21002c",
		16#42c6# => X"a9720000",
		16#42c7# => X"8521fffc",
		16#42c8# => X"8441ffd4",
		16#42c9# => X"85c1ffd8",
		16#42ca# => X"8601ffdc",
		16#42cb# => X"8641ffe0",
		16#42cc# => X"8681ffe4",
		16#42cd# => X"86c1ffe8",
		16#42ce# => X"8701ffec",
		16#42cf# => X"8741fff0",
		16#42d0# => X"8781fff4",
		16#42d1# => X"44004800",
		16#42d2# => X"87c1fff8",
		16#42d3# => X"e0885803",
		16#42d4# => X"e2c4a000",
		16#42d5# => X"e5a3b000",
		16#42d6# => X"0fffff9a",
		16#42d7# => X"15000000",
		16#42d8# => X"8467000c",
		16#42d9# => X"84870008",
		16#42da# => X"9e420008",
		16#42db# => X"d404180c",
		16#42dc# => X"03ffffdc",
		16#42dd# => X"d4032008",
		16#42de# => X"a4c60001",
		16#42df# => X"e1c67004",
		16#42e0# => X"a8a30001",
		16#42e1# => X"d4027004",
		16#42e2# => X"d4042804",
		16#42e3# => X"e0441800",
		16#42e4# => X"a8780000",
		16#42e5# => X"84a20004",
		16#42e6# => X"9c840008",
		16#42e7# => X"a8a50001",
		16#42e8# => X"07fff627",
		16#42e9# => X"d4022804",
		16#42ea# => X"03ffffd9",
		16#42eb# => X"15000000",
		16#42ec# => X"a8920000",
		16#42ed# => X"07ffdb6d",
		16#42ee# => X"a8780000",
		16#42ef# => X"bc2b0000",
		16#42f0# => X"0fffffd3",
		16#42f1# => X"aa4b0000",
		16#42f2# => X"84c20004",
		16#42f3# => X"9d80fffe",
		16#42f4# => X"9c6bfff8",
		16#42f5# => X"e0866003",
		16#42f6# => X"e0822000",
		16#42f7# => X"e4232000",
		16#42f8# => X"0c0000cd",
		16#42f9# => X"9cb4fffc",
		16#42fa# => X"bc450024",
		16#42fb# => X"1000008a",
		16#42fc# => X"a8500000",
		16#42fd# => X"bca50013",
		16#42fe# => X"10000018",
		16#42ff# => X"a86b0000",
		16#4300# => X"84500000",
		16#4301# => X"9c6b0008",
		16#4302# => X"d40b1000",
		16#4303# => X"bca5001b",
		16#4304# => X"84900004",
		16#4305# => X"9c500008",
		16#4306# => X"10000010",
		16#4307# => X"d40b2004",
		16#4308# => X"84420000",
		16#4309# => X"bc250024",
		16#430a# => X"d4031000",
		16#430b# => X"9c500010",
		16#430c# => X"8490000c",
		16#430d# => X"9c6b0010",
		16#430e# => X"10000008",
		16#430f# => X"d40b200c",
		16#4310# => X"84820000",
		16#4311# => X"9c500018",
		16#4312# => X"d4032000",
		16#4313# => X"9c6b0018",
		16#4314# => X"84900014",
		16#4315# => X"d40b2014",
		16#4316# => X"84820000",
		16#4317# => X"9c420004",
		16#4318# => X"d4032000",
		16#4319# => X"9c630004",
		16#431a# => X"84820000",
		16#431b# => X"d4032000",
		16#431c# => X"84420004",
		16#431d# => X"d4031004",
		16#431e# => X"a8780000",
		16#431f# => X"07fff5f0",
		16#4320# => X"a8900000",
		16#4321# => X"07ffdd8b",
		16#4322# => X"a8780000",
		16#4323# => X"03ffffa3",
		16#4324# => X"9c21002c",
		16#4325# => X"e3dea000",
		16#4326# => X"e543f000",
		16#4327# => X"13ffffc6",
		16#4328# => X"a8920000",
		16#4329# => X"845a000c",
		16#432a# => X"847a0008",
		16#432b# => X"9cb4fffc",
		16#432c# => X"d403100c",
		16#432d# => X"d4021808",
		16#432e# => X"bc450024",
		16#432f# => X"1000004f",
		16#4330# => X"9e5a0008",
		16#4331# => X"bca50013",
		16#4332# => X"10000018",
		16#4333# => X"a8520000",
		16#4334# => X"84700000",
		16#4335# => X"9c5a0010",
		16#4336# => X"d4121800",
		16#4337# => X"bca5001b",
		16#4338# => X"84700004",
		16#4339# => X"9e100008",
		16#433a# => X"10000010",
		16#433b# => X"d41a180c",
		16#433c# => X"84700000",
		16#433d# => X"bc250024",
		16#433e# => X"d4021800",
		16#433f# => X"9c5a0018",
		16#4340# => X"84700004",
		16#4341# => X"9e100008",
		16#4342# => X"10000008",
		16#4343# => X"d41a1814",
		16#4344# => X"84700000",
		16#4345# => X"d4021800",
		16#4346# => X"9c5a0020",
		16#4347# => X"84700004",
		16#4348# => X"9e100008",
		16#4349# => X"d41a181c",
		16#434a# => X"84700000",
		16#434b# => X"9e100004",
		16#434c# => X"d4021800",
		16#434d# => X"9c620004",
		16#434e# => X"84500000",
		16#434f# => X"aade0000",
		16#4350# => X"d4031000",
		16#4351# => X"a85a0000",
		16#4352# => X"84900004",
		16#4353# => X"d4032004",
		16#4354# => X"03ffff64",
		16#4355# => X"84da0004",
		16#4356# => X"9c21002c",
		16#4357# => X"a8850000",
		16#4358# => X"8521fffc",
		16#4359# => X"8441ffd4",
		16#435a# => X"85c1ffd8",
		16#435b# => X"8601ffdc",
		16#435c# => X"8641ffe0",
		16#435d# => X"8681ffe4",
		16#435e# => X"86c1ffe8",
		16#435f# => X"8701ffec",
		16#4360# => X"8741fff0",
		16#4361# => X"8781fff4",
		16#4362# => X"03ffdaf8",
		16#4363# => X"87c1fff8",
		16#4364# => X"9c40000c",
		16#4365# => X"9e400000",
		16#4366# => X"03ffff5f",
		16#4367# => X"d4181000",
		16#4368# => X"9ce0fffc",
		16#4369# => X"84850004",
		16#436a# => X"9d6e0010",
		16#436b# => X"e0843803",
		16#436c# => X"e104a000",
		16#436d# => X"e5885800",
		16#436e# => X"13ffff02",
		16#436f# => X"a8e50000",
		16#4370# => X"e0a87002",
		16#4371# => X"e0827000",
		16#4372# => X"a8a50001",
		16#4373# => X"d41c2008",
		16#4374# => X"d4042804",
		16#4375# => X"a8780000",
		16#4376# => X"84820004",
		16#4377# => X"aa500000",
		16#4378# => X"a4840001",
		16#4379# => X"e1ce2004",
		16#437a# => X"07ffdd32",
		16#437b# => X"d4027004",
		16#437c# => X"03ffff4a",
		16#437d# => X"9c21002c",
		16#437e# => X"a8720000",
		16#437f# => X"a8900000",
		16#4380# => X"07fff97a",
		16#4381# => X"aade0000",
		16#4382# => X"84da0004",
		16#4383# => X"03ffff35",
		16#4384# => X"a85a0000",
		16#4385# => X"a86b0000",
		16#4386# => X"07fff974",
		16#4387# => X"a8900000",
		16#4388# => X"03ffff97",
		16#4389# => X"a8780000",
		16#438a# => X"e3dea000",
		16#438b# => X"e2c4f000",
		16#438c# => X"e5962800",
		16#438d# => X"13ffff9a",
		16#438e# => X"e543f000",
		16#438f# => X"845a000c",
		16#4390# => X"847a0008",
		16#4391# => X"e0b45800",
		16#4392# => X"d403100c",
		16#4393# => X"d4021808",
		16#4394# => X"bc450024",
		16#4395# => X"1000003c",
		16#4396# => X"9e5a0008",
		16#4397# => X"bca50013",
		16#4398# => X"10000018",
		16#4399# => X"a8520000",
		16#439a# => X"84700000",
		16#439b# => X"9c5a0010",
		16#439c# => X"d4121800",
		16#439d# => X"bca5001b",
		16#439e# => X"84700004",
		16#439f# => X"9e100008",
		16#43a0# => X"10000010",
		16#43a1# => X"d41a180c",
		16#43a2# => X"84700000",
		16#43a3# => X"bc250024",
		16#43a4# => X"d4021800",
		16#43a5# => X"9c5a0018",
		16#43a6# => X"84700004",
		16#43a7# => X"9e100008",
		16#43a8# => X"10000008",
		16#43a9# => X"d41a1814",
		16#43aa# => X"84700000",
		16#43ab# => X"d4021800",
		16#43ac# => X"9c5a0020",
		16#43ad# => X"84700004",
		16#43ae# => X"9e100008",
		16#43af# => X"d41a181c",
		16#43b0# => X"84700000",
		16#43b1# => X"9e100004",
		16#43b2# => X"d4021800",
		16#43b3# => X"9c420004",
		16#43b4# => X"84700000",
		16#43b5# => X"d4021800",
		16#43b6# => X"84700004",
		16#43b7# => X"d4021804",
		16#43b8# => X"e0967002",
		16#43b9# => X"e05a7000",
		16#43ba# => X"a8840001",
		16#43bb# => X"d41c1008",
		16#43bc# => X"d4022004",
		16#43bd# => X"a8780000",
		16#43be# => X"845a0004",
		16#43bf# => X"a4420001",
		16#43c0# => X"e1ce1004",
		16#43c1# => X"07ffdceb",
		16#43c2# => X"d41a7004",
		16#43c3# => X"03ffff03",
		16#43c4# => X"9c21002c",
		16#43c5# => X"86c30004",
		16#43c6# => X"9c60fffc",
		16#43c7# => X"9e420008",
		16#43c8# => X"e2d61803",
		16#43c9# => X"03fffeef",
		16#43ca# => X"e2d6a000",
		16#43cb# => X"a8720000",
		16#43cc# => X"a8900000",
		16#43cd# => X"07fff92d",
		16#43ce# => X"a85a0000",
		16#43cf# => X"03fffee9",
		16#43d0# => X"84da0004",
		16#43d1# => X"a8720000",
		16#43d2# => X"07fff928",
		16#43d3# => X"a8900000",
		16#43d4# => X"03ffffe5",
		16#43d5# => X"e0967002",
		16#43d6# => X"d7e117f4",
		16#43d7# => X"d7e177f8",
		16#43d8# => X"d7e14ffc",
		16#43d9# => X"a8440000",
		16#43da# => X"84840000",
		16#43db# => X"9c21fff4",
		16#43dc# => X"bc040000",
		16#43dd# => X"10000004",
		16#43de# => X"a9c30000",
		16#43df# => X"07fffff7",
		16#43e0# => X"15000000",
		16#43e1# => X"9c21000c",
		16#43e2# => X"a86e0000",
		16#43e3# => X"a8820000",
		16#43e4# => X"8521fffc",
		16#43e5# => X"8441fff4",
		16#43e6# => X"03fff529",
		16#43e7# => X"85c1fff8",
		16#43e8# => X"d7e117ec",
		16#43e9# => X"18400001",
		16#43ea# => X"d7e177f0",
		16#43eb# => X"a84263e0",
		16#43ec# => X"d7e14ffc",
		16#43ed# => X"d7e187f4",
		16#43ee# => X"d7e197f8",
		16#43ef# => X"84420000",
		16#43f0# => X"9c21ffec",
		16#43f1# => X"e4031000",
		16#43f2# => X"1000003a",
		16#43f3# => X"a9c30000",
		16#43f4# => X"8483004c",
		16#43f5# => X"bc040000",
		16#43f6# => X"10000017",
		16#43f7# => X"9c400000",
		16#43f8# => X"aa020000",
		16#43f9# => X"b8420002",
		16#43fa# => X"e0441000",
		16#43fb# => X"84a20000",
		16#43fc# => X"bc050000",
		16#43fd# => X"1000000a",
		16#43fe# => X"15000000",
		16#43ff# => X"a8850000",
		16#4400# => X"a86e0000",
		16#4401# => X"07fff50e",
		16#4402# => X"84450000",
		16#4403# => X"bc220000",
		16#4404# => X"13fffffb",
		16#4405# => X"a8a20000",
		16#4406# => X"848e004c",
		16#4407# => X"9e100001",
		16#4408# => X"bc100020",
		16#4409# => X"0ffffff0",
		16#440a# => X"a8500000",
		16#440b# => X"07fff504",
		16#440c# => X"a86e0000",
		16#440d# => X"848e0040",
		16#440e# => X"bc040000",
		16#440f# => X"10000004",
		16#4410# => X"15000000",
		16#4411# => X"07fff4fe",
		16#4412# => X"a86e0000",
		16#4413# => X"844e0148",
		16#4414# => X"bc020000",
		16#4415# => X"1000000d",
		16#4416# => X"15000000",
		16#4417# => X"9e4e014c",
		16#4418# => X"e4029000",
		16#4419# => X"10000009",
		16#441a# => X"15000000",
		16#441b# => X"a8820000",
		16#441c# => X"a86e0000",
		16#441d# => X"07fff4f2",
		16#441e# => X"86020000",
		16#441f# => X"e4328000",
		16#4420# => X"13fffffb",
		16#4421# => X"a8500000",
		16#4422# => X"848e0054",
		16#4423# => X"bc040000",
		16#4424# => X"10000004",
		16#4425# => X"15000000",
		16#4426# => X"07fff4e9",
		16#4427# => X"a86e0000",
		16#4428# => X"844e0038",
		16#4429# => X"bc020000",
		16#442a# => X"0c000009",
		16#442b# => X"15000000",
		16#442c# => X"9c210014",
		16#442d# => X"8521fffc",
		16#442e# => X"8441ffec",
		16#442f# => X"85c1fff0",
		16#4430# => X"8601fff4",
		16#4431# => X"44004800",
		16#4432# => X"8641fff8",
		16#4433# => X"844e003c",
		16#4434# => X"48001000",
		16#4435# => X"a86e0000",
		16#4436# => X"848e02e0",
		16#4437# => X"bc040000",
		16#4438# => X"13fffff4",
		16#4439# => X"15000000",
		16#443a# => X"9c210014",
		16#443b# => X"a86e0000",
		16#443c# => X"8521fffc",
		16#443d# => X"8441ffec",
		16#443e# => X"85c1fff0",
		16#443f# => X"8601fff4",
		16#4440# => X"03ffff96",
		16#4441# => X"8641fff8",
		16#4442# => X"d7e197f8",
		16#4443# => X"d7e14ffc",
		16#4444# => X"d7e117ec",
		16#4445# => X"d7e177f0",
		16#4446# => X"d7e187f4",
		16#4447# => X"aa430000",
		16#4448# => X"bc230000",
		16#4449# => X"0c000029",
		16#444a# => X"9c21ffec",
		16#444b# => X"86120148",
		16#444c# => X"bc100000",
		16#444d# => X"10000013",
		16#444e# => X"15000000",
		16#444f# => X"84500004",
		16#4450# => X"9dc2ffff",
		16#4451# => X"bd8e0000",
		16#4452# => X"1000000a",
		16#4453# => X"9c420001",
		16#4454# => X"b8420002",
		16#4455# => X"e0501000",
		16#4456# => X"84820000",
		16#4457# => X"48002000",
		16#4458# => X"9dceffff",
		16#4459# => X"bd6e0000",
		16#445a# => X"13fffffc",
		16#445b# => X"9c42fffc",
		16#445c# => X"86100000",
		16#445d# => X"bc300000",
		16#445e# => X"13fffff1",
		16#445f# => X"15000000",
		16#4460# => X"8452003c",
		16#4461# => X"bc020000",
		16#4462# => X"10000009",
		16#4463# => X"a8720000",
		16#4464# => X"9c210014",
		16#4465# => X"8521fffc",
		16#4466# => X"85c1fff0",
		16#4467# => X"8601fff4",
		16#4468# => X"8641fff8",
		16#4469# => X"44001000",
		16#446a# => X"8441ffec",
		16#446b# => X"9c210014",
		16#446c# => X"8521fffc",
		16#446d# => X"8441ffec",
		16#446e# => X"85c1fff0",
		16#446f# => X"8601fff4",
		16#4470# => X"44004800",
		16#4471# => X"8641fff8",
		16#4472# => X"18400001",
		16#4473# => X"a84263e0",
		16#4474# => X"03ffffd7",
		16#4475# => X"86420000",
		16#4476# => X"d7e117fc",
		16#4477# => X"e0a41804",
		16#4478# => X"9c21fffc",
		16#4479# => X"bc050000",
		16#447a# => X"10000041",
		16#447b# => X"9d600002",
		16#447c# => X"e0a02002",
		16#447d# => X"e0852004",
		16#447e# => X"ac84ffff",
		16#447f# => X"b884005f",
		16#4480# => X"bc040000",
		16#4481# => X"0c00003d",
		16#4482# => X"18408000",
		16#4483# => X"18407ff0",
		16#4484# => X"e0c31000",
		16#4485# => X"18407fdf",
		16#4486# => X"a842ffff",
		16#4487# => X"e4a61000",
		16#4488# => X"10000003",
		16#4489# => X"9ca00001",
		16#448a# => X"9ca00000",
		16#448b# => X"a4a500ff",
		16#448c# => X"bc250000",
		16#448d# => X"10000046",
		16#448e# => X"15000000",
		16#448f# => X"1840fff0",
		16#4490# => X"e0e31000",
		16#4491# => X"18407fdf",
		16#4492# => X"a842ffff",
		16#4493# => X"e4a71000",
		16#4494# => X"0c000039",
		16#4495# => X"9cc00001",
		16#4496# => X"a4c600ff",
		16#4497# => X"bc260000",
		16#4498# => X"1000003b",
		16#4499# => X"15000000",
		16#449a# => X"18408000",
		16#449b# => X"e0e31000",
		16#449c# => X"1840000f",
		16#449d# => X"a842ffff",
		16#449e# => X"e4a71000",
		16#449f# => X"0c000027",
		16#44a0# => X"9ca00001",
		16#44a1# => X"a4a500ff",
		16#44a2# => X"bc250000",
		16#44a3# => X"1000002c",
		16#44a4# => X"15000000",
		16#44a5# => X"1840000f",
		16#44a6# => X"a842ffff",
		16#44a7# => X"e4a31000",
		16#44a8# => X"10000003",
		16#44a9# => X"9cc00001",
		16#44aa# => X"a8c50000",
		16#44ab# => X"a4c600ff",
		16#44ac# => X"bc260000",
		16#44ad# => X"10000022",
		16#44ae# => X"15000000",
		16#44af# => X"1840fff0",
		16#44b0# => X"e0a31005",
		16#44b1# => X"18407ff0",
		16#44b2# => X"e1602802",
		16#44b3# => X"e0631005",
		16#44b4# => X"e0ab2804",
		16#44b5# => X"e0c01802",
		16#44b6# => X"e0661804",
		16#44b7# => X"e1632803",
		16#44b8# => X"ad6bffff",
		16#44b9# => X"b96b005f",
		16#44ba# => X"e1645803",
		16#44bb# => X"9c210004",
		16#44bc# => X"44004800",
		16#44bd# => X"8441fffc",
		16#44be# => X"e0a31000",
		16#44bf# => X"e0c02802",
		16#44c0# => X"e0a62804",
		16#44c1# => X"bd650000",
		16#44c2# => X"0fffffc1",
		16#44c3# => X"15000000",
		16#44c4# => X"03fffff8",
		16#44c5# => X"9c210004",
		16#44c6# => X"a8a60000",
		16#44c7# => X"a4a500ff",
		16#44c8# => X"bc250000",
		16#44c9# => X"0fffffdc",
		16#44ca# => X"15000000",
		16#44cb# => X"00000005",
		16#44cc# => X"9c210004",
		16#44cd# => X"03ffffc9",
		16#44ce# => X"a8c50000",
		16#44cf# => X"9c210004",
		16#44d0# => X"9d600003",
		16#44d1# => X"44004800",
		16#44d2# => X"8441fffc",
		16#44d3# => X"9c210004",
		16#44d4# => X"9d600004",
		16#44d5# => X"44004800",
		16#44d6# => X"8441fffc",
		16#44d7# => X"d7e117f8",
		16#44d8# => X"a8440000",
		16#44d9# => X"9884000e",
		16#44da# => X"d7e14ffc",
		16#44db# => X"0400068f",
		16#44dc# => X"9c21fff8",
		16#44dd# => X"bd8b0000",
		16#44de# => X"10000009",
		16#44df# => X"9c80efff",
		16#44e0# => X"84620050",
		16#44e1# => X"e0635800",
		16#44e2# => X"d4021850",
		16#44e3# => X"9c210008",
		16#44e4# => X"8521fffc",
		16#44e5# => X"44004800",
		16#44e6# => X"8441fff8",
		16#44e7# => X"9462000c",
		16#44e8# => X"e0632003",
		16#44e9# => X"dc02180c",
		16#44ea# => X"9c210008",
		16#44eb# => X"8521fffc",
		16#44ec# => X"44004800",
		16#44ed# => X"8441fff8",
		16#44ee# => X"44004800",
		16#44ef# => X"9d600000",
		16#44f0# => X"d7e117ec",
		16#44f1# => X"a8440000",
		16#44f2# => X"9884000c",
		16#44f3# => X"d7e177f0",
		16#44f4# => X"d7e187f4",
		16#44f5# => X"d7e197f8",
		16#44f6# => X"d7e14ffc",
		16#44f7# => X"a4e40100",
		16#44f8# => X"9c21ffec",
		16#44f9# => X"aa430000",
		16#44fa# => X"aa050000",
		16#44fb# => X"bc070000",
		16#44fc# => X"10000007",
		16#44fd# => X"a9c60000",
		16#44fe# => X"9882000e",
		16#44ff# => X"9ca00000",
		16#4500# => X"0400064b",
		16#4501# => X"9cc00002",
		16#4502# => X"9882000c",
		16#4503# => X"9ca0efff",
		16#4504# => X"a8ce0000",
		16#4505# => X"e0642803",
		16#4506# => X"9882000e",
		16#4507# => X"dc02180c",
		16#4508# => X"9c210014",
		16#4509# => X"a8720000",
		16#450a# => X"a8b00000",
		16#450b# => X"8521fffc",
		16#450c# => X"8441ffec",
		16#450d# => X"85c1fff0",
		16#450e# => X"8601fff4",
		16#450f# => X"000004a9",
		16#4510# => X"8641fff8",
		16#4511# => X"d7e117f8",
		16#4512# => X"a8440000",
		16#4513# => X"9884000e",
		16#4514# => X"d7e14ffc",
		16#4515# => X"04000636",
		16#4516# => X"9c21fff8",
		16#4517# => X"bc2bffff",
		16#4518# => X"0c00000a",
		16#4519# => X"9c80efff",
		16#451a# => X"9462000c",
		16#451b# => X"a8631000",
		16#451c# => X"d4025850",
		16#451d# => X"dc02180c",
		16#451e# => X"9c210008",
		16#451f# => X"8521fffc",
		16#4520# => X"44004800",
		16#4521# => X"8441fff8",
		16#4522# => X"9462000c",
		16#4523# => X"e0632003",
		16#4524# => X"dc02180c",
		16#4525# => X"9c210008",
		16#4526# => X"8521fffc",
		16#4527# => X"44004800",
		16#4528# => X"8441fff8",
		16#4529# => X"d7e14ffc",
		16#452a# => X"9c21fffc",
		16#452b# => X"9884000e",
		16#452c# => X"9c210004",
		16#452d# => X"8521fffc",
		16#452e# => X"000004da",
		16#452f# => X"15000000",
		16#4530# => X"e1641804",
		16#4531# => X"d7e117fc",
		16#4532# => X"a56b0003",
		16#4533# => X"bc2b0000",
		16#4534# => X"10000024",
		16#4535# => X"9c21fffc",
		16#4536# => X"84a30000",
		16#4537# => X"84c40000",
		16#4538# => X"e4253000",
		16#4539# => X"1000001f",
		16#453a# => X"1840fefe",
		16#453b# => X"a842feff",
		16#453c# => X"e0c51000",
		16#453d# => X"aca5ffff",
		16#453e# => X"18408080",
		16#453f# => X"e0a62803",
		16#4540# => X"a8428080",
		16#4541# => X"e0a51003",
		16#4542# => X"bc250000",
		16#4543# => X"0c00000b",
		16#4544# => X"9c630004",
		16#4545# => X"9c63fffc",
		16#4546# => X"0000002a",
		16#4547# => X"9c210004",
		16#4548# => X"18408080",
		16#4549# => X"a8428080",
		16#454a# => X"e0c61003",
		16#454b# => X"bc260000",
		16#454c# => X"10000026",
		16#454d# => X"9c630004",
		16#454e# => X"1840fefe",
		16#454f# => X"84a30000",
		16#4550# => X"9c840004",
		16#4551# => X"a842feff",
		16#4552# => X"85040000",
		16#4553# => X"e0e51000",
		16#4554# => X"acc5ffff",
		16#4555# => X"e4054000",
		16#4556# => X"13fffff2",
		16#4557# => X"e0c73003",
		16#4558# => X"90a30000",
		16#4559# => X"bc050000",
		16#455a# => X"10000012",
		16#455b# => X"15000000",
		16#455c# => X"90c40000",
		16#455d# => X"e4262800",
		16#455e# => X"0c00000a",
		16#455f# => X"9c630001",
		16#4560# => X"9c63ffff",
		16#4561# => X"0000000c",
		16#4562# => X"8d630000",
		16#4563# => X"90c40000",
		16#4564# => X"e4062800",
		16#4565# => X"0c000007",
		16#4566# => X"15000000",
		16#4567# => X"9c630001",
		16#4568# => X"90a30000",
		16#4569# => X"bc050000",
		16#456a# => X"0ffffff9",
		16#456b# => X"9c840001",
		16#456c# => X"8d630000",
		16#456d# => X"8c640000",
		16#456e# => X"e16b1802",
		16#456f# => X"9c210004",
		16#4570# => X"44004800",
		16#4571# => X"8441fffc",
		16#4572# => X"9c210004",
		16#4573# => X"9d600000",
		16#4574# => X"44004800",
		16#4575# => X"8441fffc",
		16#4576# => X"d7e197ec",
		16#4577# => X"d7e1a7f0",
		16#4578# => X"d7e1b7f4",
		16#4579# => X"d7e14ffc",
		16#457a# => X"d7e117e0",
		16#457b# => X"d7e177e4",
		16#457c# => X"d7e187e8",
		16#457d# => X"d7e1c7f8",
		16#457e# => X"85650008",
		16#457f# => X"9c21ffe0",
		16#4580# => X"aac50000",
		16#4581# => X"aa830000",
		16#4582# => X"bc2b0000",
		16#4583# => X"0c00002f",
		16#4584# => X"aa440000",
		16#4585# => X"84440064",
		16#4586# => X"a4422000",
		16#4587# => X"bc020000",
		16#4588# => X"1000002c",
		16#4589# => X"15000000",
		16#458a# => X"87050000",
		16#458b# => X"86180004",
		16#458c# => X"ba100042",
		16#458d# => X"bdb00000",
		16#458e# => X"1000001d",
		16#458f# => X"84580000",
		16#4590# => X"00000005",
		16#4591# => X"9dc00000",
		16#4592# => X"e5507000",
		16#4593# => X"0c000017",
		16#4594# => X"15000000",
		16#4595# => X"84820000",
		16#4596# => X"a8740000",
		16#4597# => X"a8b20000",
		16#4598# => X"040004eb",
		16#4599# => X"9dce0001",
		16#459a# => X"bc0bffff",
		16#459b# => X"0ffffff7",
		16#459c# => X"9c420004",
		16#459d# => X"9c400000",
		16#459e# => X"d4161008",
		16#459f# => X"d4161004",
		16#45a0# => X"9c210020",
		16#45a1# => X"8521fffc",
		16#45a2# => X"8441ffe0",
		16#45a3# => X"85c1ffe4",
		16#45a4# => X"8601ffe8",
		16#45a5# => X"8641ffec",
		16#45a6# => X"8681fff0",
		16#45a7# => X"86c1fff4",
		16#45a8# => X"44004800",
		16#45a9# => X"8701fff8",
		16#45aa# => X"85760008",
		16#45ab# => X"ba100002",
		16#45ac# => X"e16b8002",
		16#45ad# => X"bc0b0000",
		16#45ae# => X"13ffffef",
		16#45af# => X"d4165808",
		16#45b0# => X"03ffffdb",
		16#45b1# => X"9f180008",
		16#45b2# => X"03ffffee",
		16#45b3# => X"d4055804",
		16#45b4# => X"07fff427",
		16#45b5# => X"9c400000",
		16#45b6# => X"03ffffe9",
		16#45b7# => X"d4161008",
		16#45b8# => X"d7e177d8",
		16#45b9# => X"d7e14ffc",
		16#45ba# => X"d7e117d4",
		16#45bb# => X"d7e187dc",
		16#45bc# => X"d7e197e0",
		16#45bd# => X"d7e1a7e4",
		16#45be# => X"d7e1b7e8",
		16#45bf# => X"d7e1c7ec",
		16#45c0# => X"d7e1d7f0",
		16#45c1# => X"d7e1e7f4",
		16#45c2# => X"d7e1f7f8",
		16#45c3# => X"9c21fac4",
		16#45c4# => X"a9c50000",
		16#45c5# => X"d4011824",
		16#45c6# => X"d4012020",
		16#45c7# => X"bc030000",
		16#45c8# => X"10000006",
		16#45c9# => X"d4013014",
		16#45ca# => X"84430038",
		16#45cb# => X"bc220000",
		16#45cc# => X"0c000335",
		16#45cd# => X"15000000",
		16#45ce# => X"84610020",
		16#45cf# => X"9843000c",
		16#45d0# => X"a4e2ffff",
		16#45d1# => X"a4a72000",
		16#45d2# => X"bc250000",
		16#45d3# => X"1000000b",
		16#45d4# => X"a4a70008",
		16#45d5# => X"84a30064",
		16#45d6# => X"9c60dfff",
		16#45d7# => X"a8422000",
		16#45d8# => X"84810020",
		16#45d9# => X"e0a51803",
		16#45da# => X"dc04100c",
		16#45db# => X"d4042864",
		16#45dc# => X"a4e2ffff",
		16#45dd# => X"a4a70008",
		16#45de# => X"bc050000",
		16#45df# => X"100003b1",
		16#45e0# => X"84810020",
		16#45e1# => X"84a40010",
		16#45e2# => X"bc250000",
		16#45e3# => X"0c0003ae",
		16#45e4# => X"84610024",
		16#45e5# => X"a4e7001a",
		16#45e6# => X"bc27000a",
		16#45e7# => X"0c0002ed",
		16#45e8# => X"84610020",
		16#45e9# => X"9c400000",
		16#45ea# => X"9c610500",
		16#45eb# => X"9c8104ff",
		16#45ec# => X"d4011804",
		16#45ed# => X"d4011028",
		16#45ee# => X"9c600000",
		16#45ef# => X"9c410498",
		16#45f0# => X"d4012000",
		16#45f1# => X"d4011500",
		16#45f2# => X"d4011d08",
		16#45f3# => X"d4011d04",
		16#45f4# => X"d401180c",
		16#45f5# => X"aa420000",
		16#45f6# => X"84610000",
		16#45f7# => X"84410004",
		16#45f8# => X"aace0000",
		16#45f9# => X"e0421802",
		16#45fa# => X"87410024",
		16#45fb# => X"d401102c",
		16#45fc# => X"87810020",
		16#45fd# => X"90560000",
		16#45fe# => X"aca20025",
		16#45ff# => X"a4a500ff",
		16#4600# => X"bc050000",
		16#4601# => X"10000238",
		16#4602# => X"15000000",
		16#4603# => X"a44200ff",
		16#4604# => X"bc020000",
		16#4605# => X"10000234",
		16#4606# => X"15000000",
		16#4607# => X"00000005",
		16#4608# => X"a8560000",
		16#4609# => X"bc230000",
		16#460a# => X"0c00000a",
		16#460b# => X"e1c2b002",
		16#460c# => X"9c420001",
		16#460d# => X"90a20000",
		16#460e# => X"ac650025",
		16#460f# => X"a46300ff",
		16#4610# => X"bc030000",
		16#4611# => X"0ffffff8",
		16#4612# => X"a46500ff",
		16#4613# => X"e1c2b002",
		16#4614# => X"bc0e0000",
		16#4615# => X"10000012",
		16#4616# => X"bc050000",
		16#4617# => X"84a10508",
		16#4618# => X"84c10504",
		16#4619# => X"e0a57000",
		16#461a# => X"9cc60001",
		16#461b# => X"d412b000",
		16#461c# => X"d4127004",
		16#461d# => X"d4012d08",
		16#461e# => X"bd460007",
		16#461f# => X"1000028b",
		16#4620# => X"d4013504",
		16#4621# => X"9e520008",
		16#4622# => X"8481000c",
		16#4623# => X"e0847000",
		16#4624# => X"d401200c",
		16#4625# => X"90a20000",
		16#4626# => X"bc050000",
		16#4627# => X"1000021f",
		16#4628# => X"9ca00000",
		16#4629# => X"9ec20001",
		16#462a# => X"9c400000",
		16#462b# => X"9dc0ffff",
		16#462c# => X"d801150f",
		16#462d# => X"d4012810",
		16#462e# => X"ab050000",
		16#462f# => X"90d60000",
		16#4630# => X"9ed60001",
		16#4631# => X"9c46ffe0",
		16#4632# => X"bc420058",
		16#4633# => X"0c00004d",
		16#4634# => X"18600001",
		16#4635# => X"bc060000",
		16#4636# => X"10000210",
		16#4637# => X"d8012d0f",
		16#4638# => X"9c600001",
		16#4639# => X"9c800000",
		16#463a# => X"d4011808",
		16#463b# => X"d80134d8",
		16#463c# => X"d801250f",
		16#463d# => X"abc30000",
		16#463e# => X"9e0104d8",
		16#463f# => X"9c400000",
		16#4640# => X"d4011018",
		16#4641# => X"a4580002",
		16#4642# => X"bc020000",
		16#4643# => X"10000005",
		16#4644# => X"a4980084",
		16#4645# => X"84610008",
		16#4646# => X"9c630002",
		16#4647# => X"d4011808",
		16#4648# => X"bc040000",
		16#4649# => X"0c00014c",
		16#464a# => X"d401201c",
		16#464b# => X"84610010",
		16#464c# => X"84810008",
		16#464d# => X"e2832002",
		16#464e# => X"bd540000",
		16#464f# => X"0c000146",
		16#4650# => X"bd540010",
		16#4651# => X"0c000332",
		16#4652# => X"15000000",
		16#4653# => X"19c00001",
		16#4654# => X"84a10508",
		16#4655# => X"84c10504",
		16#4656# => X"00000007",
		16#4657# => X"a9ce43b0",
		16#4658# => X"9e520008",
		16#4659# => X"9e94fff0",
		16#465a# => X"bd540010",
		16#465b# => X"0c00001a",
		16#465c# => X"9d920008",
		16#465d# => X"18600001",
		16#465e# => X"9cc60001",
		16#465f# => X"9ca50010",
		16#4660# => X"a86343b0",
		16#4661# => X"9c800010",
		16#4662# => X"d4121800",
		16#4663# => X"d4122004",
		16#4664# => X"d4012d08",
		16#4665# => X"bd460007",
		16#4666# => X"0ffffff2",
		16#4667# => X"d4013504",
		16#4668# => X"a87a0000",
		16#4669# => X"a89c0000",
		16#466a# => X"07ffff0c",
		16#466b# => X"9ca10500",
		16#466c# => X"bc2b0000",
		16#466d# => X"100001e1",
		16#466e# => X"9e94fff0",
		16#466f# => X"9d8104a0",
		16#4670# => X"9e410498",
		16#4671# => X"84a10508",
		16#4672# => X"bd540010",
		16#4673# => X"13ffffea",
		16#4674# => X"84c10504",
		16#4675# => X"9cc60001",
		16#4676# => X"e0a5a000",
		16#4677# => X"d4127000",
		16#4678# => X"d412a004",
		16#4679# => X"d4012d08",
		16#467a# => X"bd460007",
		16#467b# => X"100002b9",
		16#467c# => X"d4013504",
		16#467d# => X"9dac0008",
		16#467e# => X"0000011a",
		16#467f# => X"aa4c0000",
		16#4680# => X"b8420002",
		16#4681# => X"a863423c",
		16#4682# => X"e0421800",
		16#4683# => X"84420000",
		16#4684# => X"44001000",
		16#4685# => X"15000000",
		16#4686# => X"03ffffa9",
		16#4687# => X"ab180010",
		16#4688# => X"ab180010",
		16#4689# => X"a4b80010",
		16#468a# => X"bc050000",
		16#468b# => X"1000029e",
		16#468c# => X"a5180040",
		16#468d# => X"84610014",
		16#468e# => X"9ca00000",
		16#468f# => X"84430000",
		16#4690# => X"e1001002",
		16#4691# => X"9c630004",
		16#4692# => X"e1081004",
		16#4693# => X"d4011814",
		16#4694# => X"b908005f",
		16#4695# => X"9c600000",
		16#4696# => X"d8011d0f",
		16#4697# => X"bd8e0000",
		16#4698# => X"10000003",
		16#4699# => X"9c80ff7f",
		16#469a# => X"e3182003",
		16#469b# => X"e0c07002",
		16#469c# => X"e0c67004",
		16#469d# => X"bd860000",
		16#469e# => X"10000006",
		16#469f# => X"bc050001",
		16#46a0# => X"bc080000",
		16#46a1# => X"1000019b",
		16#46a2# => X"bc250000",
		16#46a3# => X"bc050001",
		16#46a4# => X"10000270",
		16#46a5# => X"bc050002",
		16#46a6# => X"10000262",
		16#46a7# => X"9e010500",
		16#46a8# => X"a4a20007",
		16#46a9# => X"9e10ffff",
		16#46aa# => X"9ca50030",
		16#46ab# => X"b8420043",
		16#46ac# => X"bc220000",
		16#46ad# => X"13fffffb",
		16#46ae# => X"d8102800",
		16#46af# => X"a4580001",
		16#46b0# => X"bc220000",
		16#46b1# => X"0c000008",
		16#46b2# => X"84410004",
		16#46b3# => X"bc250030",
		16#46b4# => X"0c0002d5",
		16#46b5# => X"9c800030",
		16#46b6# => X"9e10ffff",
		16#46b7# => X"d8102000",
		16#46b8# => X"84410004",
		16#46b9# => X"e3c28002",
		16#46ba# => X"d4017018",
		16#46bb# => X"84810018",
		16#46bc# => X"e57e2000",
		16#46bd# => X"10000003",
		16#46be# => X"d401f008",
		16#46bf# => X"d4012008",
		16#46c0# => X"90c1050f",
		16#46c1# => X"bc060000",
		16#46c2# => X"13ffff7f",
		16#46c3# => X"84410008",
		16#46c4# => X"9c420001",
		16#46c5# => X"03ffff7c",
		16#46c6# => X"d4011008",
		16#46c7# => X"ab180010",
		16#46c8# => X"a4580010",
		16#46c9# => X"bc020000",
		16#46ca# => X"0c000009",
		16#46cb# => X"84610014",
		16#46cc# => X"a4580040",
		16#46cd# => X"bc020000",
		16#46ce# => X"10000005",
		16#46cf# => X"84810014",
		16#46d0# => X"9ca00001",
		16#46d1# => X"0000025d",
		16#46d2# => X"84440000",
		16#46d3# => X"9ca00001",
		16#46d4# => X"03ffffbc",
		16#46d5# => X"84430000",
		16#46d6# => X"84410014",
		16#46d7# => X"84610014",
		16#46d8# => X"84420000",
		16#46d9# => X"9c630004",
		16#46da# => X"d4011010",
		16#46db# => X"bd620000",
		16#46dc# => X"13ffff53",
		16#46dd# => X"d4011814",
		16#46de# => X"e0401002",
		16#46df# => X"d4011010",
		16#46e0# => X"03ffff4f",
		16#46e1# => X"ab180004",
		16#46e2# => X"03ffff4d",
		16#46e3# => X"9ca0002b",
		16#46e4# => X"03ffff4b",
		16#46e5# => X"ab180080",
		16#46e6# => X"90d60000",
		16#46e7# => X"bc06002a",
		16#46e8# => X"100002ba",
		16#46e9# => X"9ed60001",
		16#46ea# => X"9c46ffd0",
		16#46eb# => X"bca20009",
		16#46ec# => X"0c00000b",
		16#46ed# => X"9dc00000",
		16#46ee# => X"b88e0003",
		16#46ef# => X"e1ce7000",
		16#46f0# => X"90d60000",
		16#46f1# => X"e1ce2000",
		16#46f2# => X"e1ce1000",
		16#46f3# => X"9c46ffd0",
		16#46f4# => X"bca20009",
		16#46f5# => X"13fffff9",
		16#46f6# => X"9ed60001",
		16#46f7# => X"bd6e0000",
		16#46f8# => X"13ffff3a",
		16#46f9# => X"9c46ffe0",
		16#46fa# => X"03ffff38",
		16#46fb# => X"9dc0ffff",
		16#46fc# => X"a4580010",
		16#46fd# => X"bc020000",
		16#46fe# => X"0c00024a",
		16#46ff# => X"d8012d0f",
		16#4700# => X"a4580040",
		16#4701# => X"bc020000",
		16#4702# => X"10000247",
		16#4703# => X"84610014",
		16#4704# => X"8481000c",
		16#4705# => X"84430000",
		16#4706# => X"9c630004",
		16#4707# => X"d4011814",
		16#4708# => X"03fffef5",
		16#4709# => X"dc022000",
		16#470a# => X"18800001",
		16#470b# => X"d8012d0f",
		16#470c# => X"a8843ec7",
		16#470d# => X"d4012028",
		16#470e# => X"a4580010",
		16#470f# => X"bc020000",
		16#4710# => X"0c000007",
		16#4711# => X"84610014",
		16#4712# => X"a4580040",
		16#4713# => X"bc020000",
		16#4714# => X"0c00023e",
		16#4715# => X"84810014",
		16#4716# => X"84610014",
		16#4717# => X"84430000",
		16#4718# => X"9c630004",
		16#4719# => X"d4011814",
		16#471a# => X"e1001002",
		16#471b# => X"e1081004",
		16#471c# => X"b908005f",
		16#471d# => X"bc080000",
		16#471e# => X"13ffff77",
		16#471f# => X"9ca00002",
		16#4720# => X"a4b80001",
		16#4721# => X"bc050000",
		16#4722# => X"10000008",
		16#4723# => X"9c800030",
		16#4724# => X"d801350d",
		16#4725# => X"d801250c",
		16#4726# => X"ab180002",
		16#4727# => X"9d000001",
		16#4728# => X"03ffff6d",
		16#4729# => X"9ca00002",
		16#472a# => X"03ffff6b",
		16#472b# => X"9ca00002",
		16#472c# => X"84810014",
		16#472d# => X"9c600030",
		16#472e# => X"84440000",
		16#472f# => X"9c800078",
		16#4730# => X"e1001002",
		16#4731# => X"d8011d0c",
		16#4732# => X"d801250d",
		16#4733# => X"84610014",
		16#4734# => X"18800001",
		16#4735# => X"e1081004",
		16#4736# => X"9c630004",
		16#4737# => X"a8843ec7",
		16#4738# => X"ab180002",
		16#4739# => X"b908005f",
		16#473a# => X"d4011814",
		16#473b# => X"d4012028",
		16#473c# => X"03ffff59",
		16#473d# => X"9ca00002",
		16#473e# => X"84410014",
		16#473f# => X"9c600000",
		16#4740# => X"9c820004",
		16#4741# => X"d8011d0f",
		16#4742# => X"d4012014",
		16#4743# => X"86020000",
		16#4744# => X"bc300000",
		16#4745# => X"0c000233",
		16#4746# => X"bd8e0000",
		16#4747# => X"1000022c",
		16#4748# => X"a8700000",
		16#4749# => X"9c800000",
		16#474a# => X"07fff521",
		16#474b# => X"a8ae0000",
		16#474c# => X"bc0b0000",
		16#474d# => X"10000251",
		16#474e# => X"abce0000",
		16#474f# => X"e3cb8002",
		16#4750# => X"e55e7000",
		16#4751# => X"0c000220",
		16#4752# => X"9c400000",
		16#4753# => X"9c600000",
		16#4754# => X"abce0000",
		16#4755# => X"03ffff66",
		16#4756# => X"d4011818",
		16#4757# => X"03fffed8",
		16#4758# => X"ab180001",
		16#4759# => X"bc250000",
		16#475a# => X"13fffed5",
		16#475b# => X"15000000",
		16#475c# => X"03fffed3",
		16#475d# => X"9ca00020",
		16#475e# => X"03fffed1",
		16#475f# => X"ab180040",
		16#4760# => X"d8012d0f",
		16#4761# => X"a4580010",
		16#4762# => X"bc020000",
		16#4763# => X"0c000007",
		16#4764# => X"84610014",
		16#4765# => X"a4580040",
		16#4766# => X"bc020000",
		16#4767# => X"0c0001f0",
		16#4768# => X"84810014",
		16#4769# => X"84610014",
		16#476a# => X"84430000",
		16#476b# => X"9c630004",
		16#476c# => X"bd820000",
		16#476d# => X"100001ef",
		16#476e# => X"d4011814",
		16#476f# => X"e1001002",
		16#4770# => X"9ca00001",
		16#4771# => X"e1081004",
		16#4772# => X"03ffff25",
		16#4773# => X"b908005f",
		16#4774# => X"84410014",
		16#4775# => X"9c600001",
		16#4776# => X"84a20000",
		16#4777# => X"9c800000",
		16#4778# => X"9c420004",
		16#4779# => X"d4011808",
		16#477a# => X"d8012cd8",
		16#477b# => X"d801250f",
		16#477c# => X"d4011014",
		16#477d# => X"abc30000",
		16#477e# => X"03fffec1",
		16#477f# => X"9e0104d8",
		16#4780# => X"18800001",
		16#4781# => X"d8012d0f",
		16#4782# => X"a8843eb6",
		16#4783# => X"03ffff8b",
		16#4784# => X"d4012028",
		16#4785# => X"d8012d0f",
		16#4786# => X"03ffffdb",
		16#4787# => X"ab180010",
		16#4788# => X"9c600000",
		16#4789# => X"9c46ffd0",
		16#478a# => X"b8830003",
		16#478b# => X"e0631800",
		16#478c# => X"90d60000",
		16#478d# => X"e0632000",
		16#478e# => X"e0621800",
		16#478f# => X"9c46ffd0",
		16#4790# => X"bca20009",
		16#4791# => X"13fffff9",
		16#4792# => X"9ed60001",
		16#4793# => X"03fffe9e",
		16#4794# => X"d4011810",
		16#4795# => X"9db20008",
		16#4796# => X"84a10508",
		16#4797# => X"84c10504",
		16#4798# => X"9181050f",
		16#4799# => X"bc0c0000",
		16#479a# => X"1000000f",
		16#479b# => X"bc020000",
		16#479c# => X"9cc60001",
		16#479d# => X"9ca50001",
		16#479e# => X"9c61050f",
		16#479f# => X"9c800001",
		16#47a0# => X"d4121800",
		16#47a1# => X"d4122004",
		16#47a2# => X"d4012d08",
		16#47a3# => X"bd460007",
		16#47a4# => X"1000011a",
		16#47a5# => X"d4013504",
		16#47a6# => X"aa4d0000",
		16#47a7# => X"9dad0008",
		16#47a8# => X"bc020000",
		16#47a9# => X"1000000f",
		16#47aa# => X"8481001c",
		16#47ab# => X"9cc60001",
		16#47ac# => X"9ca50002",
		16#47ad# => X"9c41050c",
		16#47ae# => X"9c600002",
		16#47af# => X"d4121000",
		16#47b0# => X"d4121804",
		16#47b1# => X"d4012d08",
		16#47b2# => X"bd460007",
		16#47b3# => X"10000116",
		16#47b4# => X"d4013504",
		16#47b5# => X"aa4d0000",
		16#47b6# => X"9dad0008",
		16#47b7# => X"8481001c",
		16#47b8# => X"bc240080",
		16#47b9# => X"0c0000ab",
		16#47ba# => X"84410010",
		16#47bb# => X"84810018",
		16#47bc# => X"e1c4f002",
		16#47bd# => X"bdae0000",
		16#47be# => X"1000002e",
		16#47bf# => X"bdae0010",
		16#47c0# => X"100001ad",
		16#47c1# => X"15000000",
		16#47c2# => X"18400001",
		16#47c3# => X"00000007",
		16#47c4# => X"a84243a0",
		16#47c5# => X"9e520008",
		16#47c6# => X"9dcefff0",
		16#47c7# => X"bd4e0010",
		16#47c8# => X"0c00001a",
		16#47c9# => X"9d920008",
		16#47ca# => X"18600001",
		16#47cb# => X"9cc60001",
		16#47cc# => X"9ca50010",
		16#47cd# => X"a86343a0",
		16#47ce# => X"9c800010",
		16#47cf# => X"d4121800",
		16#47d0# => X"d4122004",
		16#47d1# => X"d4012d08",
		16#47d2# => X"bd460007",
		16#47d3# => X"0ffffff2",
		16#47d4# => X"d4013504",
		16#47d5# => X"a87a0000",
		16#47d6# => X"a89c0000",
		16#47d7# => X"07fffd9f",
		16#47d8# => X"9ca10500",
		16#47d9# => X"bc2b0000",
		16#47da# => X"10000074",
		16#47db# => X"9dcefff0",
		16#47dc# => X"9d8104a0",
		16#47dd# => X"9e410498",
		16#47de# => X"84a10508",
		16#47df# => X"bd4e0010",
		16#47e0# => X"13ffffea",
		16#47e1# => X"84c10504",
		16#47e2# => X"9cc60001",
		16#47e3# => X"e0a57000",
		16#47e4# => X"d4121000",
		16#47e5# => X"d4127004",
		16#47e6# => X"d4012d08",
		16#47e7# => X"bd460007",
		16#47e8# => X"100000cb",
		16#47e9# => X"d4013504",
		16#47ea# => X"9dac0008",
		16#47eb# => X"aa4c0000",
		16#47ec# => X"9cc60001",
		16#47ed# => X"e0a5f000",
		16#47ee# => X"d4128000",
		16#47ef# => X"d412f004",
		16#47f0# => X"d4012d08",
		16#47f1# => X"bda60007",
		16#47f2# => X"0c0000a4",
		16#47f3# => X"d4013504",
		16#47f4# => X"a4d80004",
		16#47f5# => X"bc260000",
		16#47f6# => X"0c000032",
		16#47f7# => X"84410008",
		16#47f8# => X"84610010",
		16#47f9# => X"84810008",
		16#47fa# => X"e0432002",
		16#47fb# => X"bd420000",
		16#47fc# => X"0c00002b",
		16#47fd# => X"bda20010",
		16#47fe# => X"1000018e",
		16#47ff# => X"15000000",
		16#4800# => X"19c00001",
		16#4801# => X"84c10504",
		16#4802# => X"00000006",
		16#4803# => X"a9ce43b0",
		16#4804# => X"9c42fff0",
		16#4805# => X"bd420010",
		16#4806# => X"0c000019",
		16#4807# => X"9dad0008",
		16#4808# => X"18600001",
		16#4809# => X"9cc60001",
		16#480a# => X"9ca50010",
		16#480b# => X"a86343b0",
		16#480c# => X"9c800010",
		16#480d# => X"d40d1800",
		16#480e# => X"d40d2004",
		16#480f# => X"d4012d08",
		16#4810# => X"bd460007",
		16#4811# => X"0ffffff3",
		16#4812# => X"d4013504",
		16#4813# => X"a87a0000",
		16#4814# => X"a89c0000",
		16#4815# => X"07fffd61",
		16#4816# => X"9ca10500",
		16#4817# => X"bc2b0000",
		16#4818# => X"10000036",
		16#4819# => X"9c42fff0",
		16#481a# => X"9da10498",
		16#481b# => X"84a10508",
		16#481c# => X"bd420010",
		16#481d# => X"13ffffeb",
		16#481e# => X"84c10504",
		16#481f# => X"9cc60001",
		16#4820# => X"e0a22800",
		16#4821# => X"d40d7000",
		16#4822# => X"d40d1004",
		16#4823# => X"d4012d08",
		16#4824# => X"bda60007",
		16#4825# => X"0c00011a",
		16#4826# => X"d4013504",
		16#4827# => X"84410008",
		16#4828# => X"84610010",
		16#4829# => X"e5621800",
		16#482a# => X"10000003",
		16#482b# => X"8481000c",
		16#482c# => X"a8430000",
		16#482d# => X"bc050000",
		16#482e# => X"e0841000",
		16#482f# => X"0c000070",
		16#4830# => X"d401200c",
		16#4831# => X"9c400000",
		16#4832# => X"d4011504",
		16#4833# => X"90560000",
		16#4834# => X"aca20025",
		16#4835# => X"a4a500ff",
		16#4836# => X"bc050000",
		16#4837# => X"0ffffdcc",
		16#4838# => X"9e410498",
		16#4839# => X"a8560000",
		16#483a# => X"03fffdec",
		16#483b# => X"90b60000",
		16#483c# => X"1000006c",
		16#483d# => X"abc80000",
		16#483e# => X"a4580001",
		16#483f# => X"bc020000",
		16#4840# => X"100000c5",
		16#4841# => X"9c400030",
		16#4842# => X"87c1002c",
		16#4843# => X"d80114ff",
		16#4844# => X"03fffe76",
		16#4845# => X"9e0104ff",
		16#4846# => X"84410508",
		16#4847# => X"bc020000",
		16#4848# => X"10000007",
		16#4849# => X"84610020",
		16#484a# => X"84610024",
		16#484b# => X"84810020",
		16#484c# => X"07fffd2a",
		16#484d# => X"9ca10500",
		16#484e# => X"84610020",
		16#484f# => X"9443000c",
		16#4850# => X"a4420040",
		16#4851# => X"bc020000",
		16#4852# => X"10000005",
		16#4853# => X"8561000c",
		16#4854# => X"9c80ffff",
		16#4855# => X"d401200c",
		16#4856# => X"8561000c",
		16#4857# => X"9c21053c",
		16#4858# => X"8521fffc",
		16#4859# => X"8441ffd4",
		16#485a# => X"85c1ffd8",
		16#485b# => X"8601ffdc",
		16#485c# => X"8641ffe0",
		16#485d# => X"8681ffe4",
		16#485e# => X"86c1ffe8",
		16#485f# => X"8701ffec",
		16#4860# => X"8741fff0",
		16#4861# => X"8781fff4",
		16#4862# => X"44004800",
		16#4863# => X"87c1fff8",
		16#4864# => X"84610008",
		16#4865# => X"e2821802",
		16#4866# => X"bd540000",
		16#4867# => X"0c0000f9",
		16#4868# => X"bdb40010",
		16#4869# => X"10000131",
		16#486a# => X"15000000",
		16#486b# => X"18400001",
		16#486c# => X"00000007",
		16#486d# => X"a84243a0",
		16#486e# => X"9e520008",
		16#486f# => X"9e94fff0",
		16#4870# => X"bd540010",
		16#4871# => X"0c00001a",
		16#4872# => X"9d920008",
		16#4873# => X"18800001",
		16#4874# => X"9cc60001",
		16#4875# => X"9ca50010",
		16#4876# => X"a88443a0",
		16#4877# => X"9c600010",
		16#4878# => X"d4122000",
		16#4879# => X"d4121804",
		16#487a# => X"d4012d08",
		16#487b# => X"bd460007",
		16#487c# => X"0ffffff2",
		16#487d# => X"d4013504",
		16#487e# => X"a87a0000",
		16#487f# => X"a89c0000",
		16#4880# => X"07fffcf6",
		16#4881# => X"9ca10500",
		16#4882# => X"bc2b0000",
		16#4883# => X"13ffffcb",
		16#4884# => X"9e94fff0",
		16#4885# => X"9d8104a0",
		16#4886# => X"9e410498",
		16#4887# => X"84a10508",
		16#4888# => X"bd540010",
		16#4889# => X"13ffffea",
		16#488a# => X"84c10504",
		16#488b# => X"9cc60001",
		16#488c# => X"e0a5a000",
		16#488d# => X"d4121000",
		16#488e# => X"d412a004",
		16#488f# => X"d4012d08",
		16#4890# => X"bd460007",
		16#4891# => X"100000d1",
		16#4892# => X"d4013504",
		16#4893# => X"9dac0008",
		16#4894# => X"03ffff27",
		16#4895# => X"aa4c0000",
		16#4896# => X"a87a0000",
		16#4897# => X"a89c0000",
		16#4898# => X"07fffcde",
		16#4899# => X"9ca10500",
		16#489a# => X"bc2b0000",
		16#489b# => X"13ffffb3",
		16#489c# => X"9da10498",
		16#489d# => X"03ffff57",
		16#489e# => X"84a10508",
		16#489f# => X"a87a0000",
		16#48a0# => X"a89c0000",
		16#48a1# => X"07fffcd5",
		16#48a2# => X"9ca10500",
		16#48a3# => X"bc2b0000",
		16#48a4# => X"0fffff8e",
		16#48a5# => X"9c400000",
		16#48a6# => X"03ffffa9",
		16#48a7# => X"84610020",
		16#48a8# => X"03fffe12",
		16#48a9# => X"9e010500",
		16#48aa# => X"a87a0000",
		16#48ab# => X"a89c0000",
		16#48ac# => X"07fffcca",
		16#48ad# => X"9ca10500",
		16#48ae# => X"bc2b0000",
		16#48af# => X"13ffff9f",
		16#48b0# => X"9e410498",
		16#48b1# => X"03fffd72",
		16#48b2# => X"8481000c",
		16#48b3# => X"a87a0000",
		16#48b4# => X"a89c0000",
		16#48b5# => X"07fffcc1",
		16#48b6# => X"9ca10500",
		16#48b7# => X"bc2b0000",
		16#48b8# => X"13ffff96",
		16#48b9# => X"9da104a0",
		16#48ba# => X"9e410498",
		16#48bb# => X"84a10508",
		16#48bc# => X"03ffff30",
		16#48bd# => X"84c10504",
		16#48be# => X"a87a0000",
		16#48bf# => X"a89c0000",
		16#48c0# => X"07fffcb6",
		16#48c1# => X"9ca10500",
		16#48c2# => X"bc2b0000",
		16#48c3# => X"13ffff8b",
		16#48c4# => X"9da104a0",
		16#48c5# => X"9e410498",
		16#48c6# => X"84a10508",
		16#48c7# => X"03fffee1",
		16#48c8# => X"84c10504",
		16#48c9# => X"a87a0000",
		16#48ca# => X"a89c0000",
		16#48cb# => X"07fffcab",
		16#48cc# => X"9ca10500",
		16#48cd# => X"bc2b0000",
		16#48ce# => X"13ffff80",
		16#48cf# => X"9da104a0",
		16#48d0# => X"9e410498",
		16#48d1# => X"84a10508",
		16#48d2# => X"03fffee5",
		16#48d3# => X"84c10504",
		16#48d4# => X"98e3000e",
		16#48d5# => X"bd870000",
		16#48d6# => X"13fffd13",
		16#48d7# => X"9c80fffd",
		16#48d8# => X"9e010430",
		16#48d9# => X"e0422003",
		16#48da# => X"85e30064",
		16#48db# => X"85a3001c",
		16#48dc# => X"85830024",
		16#48dd# => X"9d610030",
		16#48de# => X"9d000400",
		16#48df# => X"dc01143c",
		16#48e0# => X"84610024",
		16#48e1# => X"9c400000",
		16#48e2# => X"a8900000",
		16#48e3# => X"a8ae0000",
		16#48e4# => X"84c10014",
		16#48e5# => X"d4017c94",
		16#48e6# => X"dc013c3e",
		16#48e7# => X"d4016c4c",
		16#48e8# => X"d4016454",
		16#48e9# => X"d4015c30",
		16#48ea# => X"d4015c40",
		16#48eb# => X"d4014438",
		16#48ec# => X"d4014444",
		16#48ed# => X"07fffccb",
		16#48ee# => X"d4011448",
		16#48ef# => X"e58b1000",
		16#48f0# => X"10000008",
		16#48f1# => X"d401580c",
		16#48f2# => X"84610024",
		16#48f3# => X"07ffeded",
		16#48f4# => X"a8900000",
		16#48f5# => X"e42b1000",
		16#48f6# => X"100000aa",
		16#48f7# => X"9c60ffff",
		16#48f8# => X"9441043c",
		16#48f9# => X"a4420040",
		16#48fa# => X"bc020000",
		16#48fb# => X"13ffff5b",
		16#48fc# => X"84810020",
		16#48fd# => X"9444000c",
		16#48fe# => X"a8420040",
		16#48ff# => X"03ffff57",
		16#4900# => X"dc04100c",
		16#4901# => X"07ffeeed",
		16#4902# => X"15000000",
		16#4903# => X"03fffccc",
		16#4904# => X"84610020",
		16#4905# => X"abc50000",
		16#4906# => X"03fffdb4",
		16#4907# => X"9e010500",
		16#4908# => X"84810028",
		16#4909# => X"a462000f",
		16#490a# => X"9e10ffff",
		16#490b# => X"e0641800",
		16#490c# => X"b8420044",
		16#490d# => X"8c630000",
		16#490e# => X"bc220000",
		16#490f# => X"13fffffa",
		16#4910# => X"d8101800",
		16#4911# => X"84810004",
		16#4912# => X"03fffda8",
		16#4913# => X"e3c48002",
		16#4914# => X"bc420009",
		16#4915# => X"0c00000e",
		16#4916# => X"9e010500",
		16#4917# => X"a8620000",
		16#4918# => X"9c80000a",
		16#4919# => X"0400052d",
		16#491a# => X"9e10ffff",
		16#491b# => X"9d6b0030",
		16#491c# => X"a8620000",
		16#491d# => X"9c80000a",
		16#491e# => X"07ffc9a3",
		16#491f# => X"d8105800",
		16#4920# => X"bc4b0009",
		16#4921# => X"13fffff6",
		16#4922# => X"a84b0000",
		16#4923# => X"9e10ffff",
		16#4924# => X"84610004",
		16#4925# => X"9c420030",
		16#4926# => X"e3c38002",
		16#4927# => X"03fffd93",
		16#4928# => X"d8101000",
		16#4929# => X"bc080000",
		16#492a# => X"10000025",
		16#492b# => X"84610014",
		16#492c# => X"84810014",
		16#492d# => X"84440000",
		16#492e# => X"a442ffff",
		16#492f# => X"9c840004",
		16#4930# => X"e1001002",
		16#4931# => X"d4012014",
		16#4932# => X"03fffd63",
		16#4933# => X"b908005f",
		16#4934# => X"a87a0000",
		16#4935# => X"a89c0000",
		16#4936# => X"07fffc40",
		16#4937# => X"9ca10500",
		16#4938# => X"bc2b0000",
		16#4939# => X"13ffff15",
		16#493a# => X"9da104a0",
		16#493b# => X"9e410498",
		16#493c# => X"84a10508",
		16#493d# => X"03fffe5b",
		16#493e# => X"84c10504",
		16#493f# => X"a87a0000",
		16#4940# => X"a89c0000",
		16#4941# => X"07fffc35",
		16#4942# => X"9ca10500",
		16#4943# => X"bc2b0000",
		16#4944# => X"13ffff0b",
		16#4945# => X"84610020",
		16#4946# => X"03fffee1",
		16#4947# => X"84a10508",
		16#4948# => X"84610014",
		16#4949# => X"8481000c",
		16#494a# => X"84430000",
		16#494b# => X"9c630004",
		16#494c# => X"d4011814",
		16#494d# => X"03fffcb0",
		16#494e# => X"d4022000",
		16#494f# => X"a8a80000",
		16#4950# => X"03fffd40",
		16#4951# => X"84430000",
		16#4952# => X"84440000",
		16#4953# => X"9c840004",
		16#4954# => X"a442ffff",
		16#4955# => X"03fffdc5",
		16#4956# => X"d4012014",
		16#4957# => X"98440002",
		16#4958# => X"9c840004",
		16#4959# => X"bd820000",
		16#495a# => X"0ffffe15",
		16#495b# => X"d4012014",
		16#495c# => X"9c80002d",
		16#495d# => X"e0401002",
		16#495e# => X"03fffe11",
		16#495f# => X"d801250f",
		16#4960# => X"03fffe5b",
		16#4961# => X"9db20008",
		16#4962# => X"a87a0000",
		16#4963# => X"a89c0000",
		16#4964# => X"07fffc12",
		16#4965# => X"9ca10500",
		16#4966# => X"bc2b0000",
		16#4967# => X"13fffee7",
		16#4968# => X"9da104a0",
		16#4969# => X"9e410498",
		16#496a# => X"84a10508",
		16#496b# => X"03fffe50",
		16#496c# => X"84c10504",
		16#496d# => X"18400001",
		16#496e# => X"a98d0000",
		16#496f# => X"03fffe73",
		16#4970# => X"a84243a0",
		16#4971# => X"03fffd4a",
		16#4972# => X"d4011018",
		16#4973# => X"9c400000",
		16#4974# => X"07ffdbe9",
		16#4975# => X"d4011018",
		16#4976# => X"03fffd45",
		16#4977# => X"abcb0000",
		16#4978# => X"bcae0006",
		16#4979# => X"10000003",
		16#497a# => X"abce0000",
		16#497b# => X"9fc00006",
		16#497c# => X"ac5effff",
		16#497d# => X"1a000001",
		16#497e# => X"b842009f",
		16#497f# => X"aa103ed8",
		16#4980# => X"e05e1003",
		16#4981# => X"03fffcbe",
		16#4982# => X"d4011008",
		16#4983# => X"19c00001",
		16#4984# => X"9d920008",
		16#4985# => X"84a10508",
		16#4986# => X"84c10504",
		16#4987# => X"03fffcee",
		16#4988# => X"a9ce43b0",
		16#4989# => X"84610004",
		16#498a# => X"03fffd30",
		16#498b# => X"e3c38002",
		16#498c# => X"19c00001",
		16#498d# => X"84c10504",
		16#498e# => X"03fffe91",
		16#498f# => X"a9ce43b0",
		16#4990# => X"84610024",
		16#4991# => X"9c40ffff",
		16#4992# => X"07ffe454",
		16#4993# => X"d401100c",
		16#4994# => X"bc2b0000",
		16#4995# => X"13fffec1",
		16#4996# => X"84610020",
		16#4997# => X"9843000c",
		16#4998# => X"03fffc4d",
		16#4999# => X"a4e2ffff",
		16#499a# => X"18400001",
		16#499b# => X"a98d0000",
		16#499c# => X"03fffeef",
		16#499d# => X"a84243a0",
		16#499e# => X"03fffd1d",
		16#499f# => X"d4015818",
		16#49a0# => X"03ffff58",
		16#49a1# => X"d401180c",
		16#49a2# => X"84810014",
		16#49a3# => X"85c40000",
		16#49a4# => X"bd8e0000",
		16#49a5# => X"10000004",
		16#49a6# => X"9c440004",
		16#49a7# => X"03fffc88",
		16#49a8# => X"d4011014",
		16#49a9# => X"d4011014",
		16#49aa# => X"03fffc85",
		16#49ab# => X"9dc0ffff",
		16#49ac# => X"a8e40000",
		16#49ad# => X"a8830000",
		16#49ae# => X"18600001",
		16#49af# => X"d7e14ffc",
		16#49b0# => X"a86363e0",
		16#49b1# => X"9c21fffc",
		16#49b2# => X"84630000",
		16#49b3# => X"9c210004",
		16#49b4# => X"a8c50000",
		16#49b5# => X"8521fffc",
		16#49b6# => X"03fffc02",
		16#49b7# => X"a8a70000",
		16#49b8# => X"d7e117f4",
		16#49b9# => X"18400001",
		16#49ba# => X"d7e177f8",
		16#49bb# => X"a8429ad0",
		16#49bc# => X"a9c30000",
		16#49bd# => X"a8640000",
		16#49be# => X"a8850000",
		16#49bf# => X"a8a60000",
		16#49c0# => X"9cc00000",
		16#49c1# => X"d7e14ffc",
		16#49c2# => X"d4023000",
		16#49c3# => X"04000444",
		16#49c4# => X"9c21fff4",
		16#49c5# => X"bc2bffff",
		16#49c6# => X"0c000007",
		16#49c7# => X"15000000",
		16#49c8# => X"9c21000c",
		16#49c9# => X"8521fffc",
		16#49ca# => X"8441fff4",
		16#49cb# => X"44004800",
		16#49cc# => X"85c1fff8",
		16#49cd# => X"84420000",
		16#49ce# => X"bc020000",
		16#49cf# => X"13fffff9",
		16#49d0# => X"15000000",
		16#49d1# => X"d40e1000",
		16#49d2# => X"9c21000c",
		16#49d3# => X"8521fffc",
		16#49d4# => X"8441fff4",
		16#49d5# => X"44004800",
		16#49d6# => X"85c1fff8",
		16#49d7# => X"e0852306",
		16#49d8# => X"d7e117f8",
		16#49d9# => X"d7e14ffc",
		16#49da# => X"07ffd480",
		16#49db# => X"9c21fff8",
		16#49dc# => X"bc0b0000",
		16#49dd# => X"1000001e",
		16#49de# => X"a84b0000",
		16#49df# => X"9c60fffc",
		16#49e0# => X"84abfffc",
		16#49e1# => X"e0a51803",
		16#49e2# => X"e0a51800",
		16#49e3# => X"bc450024",
		16#49e4# => X"1000001c",
		16#49e5# => X"bca50013",
		16#49e6# => X"10000010",
		16#49e7# => X"a86b0000",
		16#49e8# => X"9c800000",
		16#49e9# => X"9c6b0008",
		16#49ea# => X"d40b2000",
		16#49eb# => X"bca5001b",
		16#49ec# => X"1000000a",
		16#49ed# => X"d40b2004",
		16#49ee# => X"d4032000",
		16#49ef# => X"d40b200c",
		16#49f0# => X"bc250024",
		16#49f1# => X"10000005",
		16#49f2# => X"9c6b0010",
		16#49f3# => X"d4032000",
		16#49f4# => X"d40b2014",
		16#49f5# => X"9c6b0018",
		16#49f6# => X"9ca00000",
		16#49f7# => X"9c830004",
		16#49f8# => X"d4032800",
		16#49f9# => X"d4042800",
		16#49fa# => X"d4042804",
		16#49fb# => X"9c210008",
		16#49fc# => X"a9620000",
		16#49fd# => X"8521fffc",
		16#49fe# => X"44004800",
		16#49ff# => X"8441fff8",
		16#4a00# => X"a86b0000",
		16#4a01# => X"07fff358",
		16#4a02# => X"9c800000",
		16#4a03# => X"9c210008",
		16#4a04# => X"a9620000",
		16#4a05# => X"8521fffc",
		16#4a06# => X"44004800",
		16#4a07# => X"8441fff8",
		16#4a08# => X"d7e117f4",
		16#4a09# => X"18400001",
		16#4a0a# => X"d7e177f8",
		16#4a0b# => X"a8429ad0",
		16#4a0c# => X"a9c30000",
		16#4a0d# => X"a8640000",
		16#4a0e# => X"9c800000",
		16#4a0f# => X"d7e14ffc",
		16#4a10# => X"d4022000",
		16#4a11# => X"04000283",
		16#4a12# => X"9c21fff4",
		16#4a13# => X"bc2bffff",
		16#4a14# => X"0c000007",
		16#4a15# => X"15000000",
		16#4a16# => X"9c21000c",
		16#4a17# => X"8521fffc",
		16#4a18# => X"8441fff4",
		16#4a19# => X"44004800",
		16#4a1a# => X"85c1fff8",
		16#4a1b# => X"84420000",
		16#4a1c# => X"bc020000",
		16#4a1d# => X"13fffff9",
		16#4a1e# => X"15000000",
		16#4a1f# => X"d40e1000",
		16#4a20# => X"9c21000c",
		16#4a21# => X"8521fffc",
		16#4a22# => X"8441fff4",
		16#4a23# => X"44004800",
		16#4a24# => X"85c1fff8",
		16#4a25# => X"d7e117f0",
		16#4a26# => X"d7e177f4",
		16#4a27# => X"d7e187f8",
		16#4a28# => X"d7e14ffc",
		16#4a29# => X"a8440000",
		16#4a2a# => X"9c21fff0",
		16#4a2b# => X"a9c30000",
		16#4a2c# => X"bc040000",
		16#4a2d# => X"10000037",
		16#4a2e# => X"aa040000",
		16#4a2f# => X"07ffee74",
		16#4a30# => X"15000000",
		16#4a31# => X"bc0e0000",
		16#4a32# => X"10000006",
		16#4a33# => X"15000000",
		16#4a34# => X"846e0038",
		16#4a35# => X"bc230000",
		16#4a36# => X"0c000035",
		16#4a37# => X"15000000",
		16#4a38# => X"9a02000c",
		16#4a39# => X"bc300000",
		16#4a3a# => X"0c000028",
		16#4a3b# => X"a86e0000",
		16#4a3c# => X"07ffeca4",
		16#4a3d# => X"a8820000",
		16#4a3e# => X"aa0b0000",
		16#4a3f# => X"8562002c",
		16#4a40# => X"bc0b0000",
		16#4a41# => X"10000007",
		16#4a42# => X"a86e0000",
		16#4a43# => X"48005800",
		16#4a44# => X"8482001c",
		16#4a45# => X"bd8b0000",
		16#4a46# => X"10000031",
		16#4a47# => X"15000000",
		16#4a48# => X"9462000c",
		16#4a49# => X"a4630080",
		16#4a4a# => X"bc030000",
		16#4a4b# => X"0c000028",
		16#4a4c# => X"a86e0000",
		16#4a4d# => X"84820030",
		16#4a4e# => X"bc040000",
		16#4a4f# => X"10000009",
		16#4a50# => X"9c620040",
		16#4a51# => X"e4041800",
		16#4a52# => X"10000005",
		16#4a53# => X"9c600000",
		16#4a54# => X"07ffeebb",
		16#4a55# => X"a86e0000",
		16#4a56# => X"9c600000",
		16#4a57# => X"d4021830",
		16#4a58# => X"84820044",
		16#4a59# => X"bc040000",
		16#4a5a# => X"10000007",
		16#4a5b# => X"9c600000",
		16#4a5c# => X"07ffeeb3",
		16#4a5d# => X"a86e0000",
		16#4a5e# => X"9c600000",
		16#4a5f# => X"d4021844",
		16#4a60# => X"9c600000",
		16#4a61# => X"dc02180c",
		16#4a62# => X"07ffee43",
		16#4a63# => X"15000000",
		16#4a64# => X"9c210010",
		16#4a65# => X"a9700000",
		16#4a66# => X"8521fffc",
		16#4a67# => X"8441fff0",
		16#4a68# => X"85c1fff4",
		16#4a69# => X"44004800",
		16#4a6a# => X"8601fff8",
		16#4a6b# => X"07ffed83",
		16#4a6c# => X"a86e0000",
		16#4a6d# => X"9a02000c",
		16#4a6e# => X"bc300000",
		16#4a6f# => X"13ffffcd",
		16#4a70# => X"a86e0000",
		16#4a71# => X"03fffff1",
		16#4a72# => X"15000000",
		16#4a73# => X"07ffee9c",
		16#4a74# => X"84820010",
		16#4a75# => X"03ffffd9",
		16#4a76# => X"84820030",
		16#4a77# => X"03ffffd1",
		16#4a78# => X"9e00ffff",
		16#4a79# => X"a8830000",
		16#4a7a# => X"18600001",
		16#4a7b# => X"d7e14ffc",
		16#4a7c# => X"a86363e0",
		16#4a7d# => X"9c21fffc",
		16#4a7e# => X"84630000",
		16#4a7f# => X"9c210004",
		16#4a80# => X"8521fffc",
		16#4a81# => X"03ffffa4",
		16#4a82# => X"15000000",
		16#4a83# => X"d7e1b7f8",
		16#4a84# => X"aac30000",
		16#4a85# => X"9865000c",
		16#4a86# => X"d7e117e4",
		16#4a87# => X"d7e1a7f4",
		16#4a88# => X"d7e14ffc",
		16#4a89# => X"d7e177e8",
		16#4a8a# => X"d7e187ec",
		16#4a8b# => X"d7e197f0",
		16#4a8c# => X"a8450000",
		16#4a8d# => X"a4a32000",
		16#4a8e# => X"9c21ffe0",
		16#4a8f# => X"bc250000",
		16#4a90# => X"10000007",
		16#4a91# => X"aa840000",
		16#4a92# => X"84820064",
		16#4a93# => X"a8632000",
		16#4a94# => X"a8842000",
		16#4a95# => X"dc02180c",
		16#4a96# => X"d4022064",
		16#4a97# => X"bdb40000",
		16#4a98# => X"1000003e",
		16#4a99# => X"18600001",
		16#4a9a# => X"a8636d90",
		16#4a9b# => X"84630000",
		16#4a9c# => X"ac630001",
		16#4a9d# => X"e0801802",
		16#4a9e# => X"e0641804",
		16#4a9f# => X"bd830000",
		16#4aa0# => X"10000036",
		16#4aa1# => X"bd5400ff",
		16#4aa2# => X"10000034",
		16#4aa3# => X"9e400001",
		16#4aa4# => X"d801a003",
		16#4aa5# => X"9dc10003",
		16#4aa6# => X"0000000c",
		16#4aa7# => X"9e000000",
		16#4aa8# => X"8c6e0000",
		16#4aa9# => X"84820000",
		16#4aaa# => X"d8041800",
		16#4aab# => X"84c20000",
		16#4aac# => X"9cc60001",
		16#4aad# => X"d4023000",
		16#4aae# => X"9e100001",
		16#4aaf# => X"e4909000",
		16#4ab0# => X"0c000032",
		16#4ab1# => X"9dce0001",
		16#4ab2# => X"84c20008",
		16#4ab3# => X"9cc6ffff",
		16#4ab4# => X"bd660000",
		16#4ab5# => X"13fffff3",
		16#4ab6# => X"d4023008",
		16#4ab7# => X"84620018",
		16#4ab8# => X"e5861800",
		16#4ab9# => X"1000002f",
		16#4aba# => X"15000000",
		16#4abb# => X"8c8e0000",
		16#4abc# => X"84620000",
		16#4abd# => X"d8032000",
		16#4abe# => X"84820000",
		16#4abf# => X"8cc40000",
		16#4ac0# => X"ac66ffff",
		16#4ac1# => X"9ca40001",
		16#4ac2# => X"e0801802",
		16#4ac3# => X"bc06000a",
		16#4ac4# => X"1000002e",
		16#4ac5# => X"e0641804",
		16#4ac6# => X"ac63ffff",
		16#4ac7# => X"d4022800",
		16#4ac8# => X"b8c3005f",
		16#4ac9# => X"bc260000",
		16#4aca# => X"0fffffe5",
		16#4acb# => X"9e100001",
		16#4acc# => X"9d60ffff",
		16#4acd# => X"9c210020",
		16#4ace# => X"8521fffc",
		16#4acf# => X"8441ffe4",
		16#4ad0# => X"85c1ffe8",
		16#4ad1# => X"8601ffec",
		16#4ad2# => X"8641fff0",
		16#4ad3# => X"8681fff4",
		16#4ad4# => X"44004800",
		16#4ad5# => X"86c1fff8",
		16#4ad6# => X"9dc10003",
		16#4ad7# => X"a8760000",
		16#4ad8# => X"a88e0000",
		16#4ad9# => X"a8b40000",
		16#4ada# => X"04000124",
		16#4adb# => X"9cc2005c",
		16#4adc# => X"bc2bffff",
		16#4add# => X"0c000007",
		16#4ade# => X"aa4b0000",
		16#4adf# => X"bc2b0000",
		16#4ae0# => X"13ffffd2",
		16#4ae1# => X"9e000000",
		16#4ae2# => X"03ffffeb",
		16#4ae3# => X"a9740000",
		16#4ae4# => X"9462000c",
		16#4ae5# => X"a8630040",
		16#4ae6# => X"03ffffe7",
		16#4ae7# => X"dc02180c",
		16#4ae8# => X"8c8e0000",
		16#4ae9# => X"a8760000",
		16#4aea# => X"0400009f",
		16#4aeb# => X"a8a20000",
		16#4aec# => X"ad6bffff",
		16#4aed# => X"e0c05802",
		16#4aee# => X"e0c65804",
		16#4aef# => X"acc6ffff",
		16#4af0# => X"03ffffd9",
		16#4af1# => X"b8c6005f",
		16#4af2# => X"a8760000",
		16#4af3# => X"03fffff7",
		16#4af4# => X"a8860000",
		16#4af5# => X"d7e187f8",
		16#4af6# => X"1a000001",
		16#4af7# => X"d7e117f0",
		16#4af8# => X"aa1063e0",
		16#4af9# => X"d7e177f4",
		16#4afa# => X"d7e14ffc",
		16#4afb# => X"a9c30000",
		16#4afc# => X"84700000",
		16#4afd# => X"9c21fff0",
		16#4afe# => X"bc030000",
		16#4aff# => X"10000009",
		16#4b00# => X"a8440000",
		16#4b01# => X"84830038",
		16#4b02# => X"bc240000",
		16#4b03# => X"10000005",
		16#4b04# => X"15000000",
		16#4b05# => X"07ffece9",
		16#4b06# => X"15000000",
		16#4b07# => X"84700000",
		16#4b08# => X"9c210010",
		16#4b09# => X"a88e0000",
		16#4b0a# => X"a8a20000",
		16#4b0b# => X"8521fffc",
		16#4b0c# => X"8441fff0",
		16#4b0d# => X"85c1fff4",
		16#4b0e# => X"03ffff75",
		16#4b0f# => X"8601fff8",
		16#4b10# => X"d7e117f4",
		16#4b11# => X"18400001",
		16#4b12# => X"d7e177f8",
		16#4b13# => X"a8429ad0",
		16#4b14# => X"a9c30000",
		16#4b15# => X"a8640000",
		16#4b16# => X"a8850000",
		16#4b17# => X"9ca00000",
		16#4b18# => X"d7e14ffc",
		16#4b19# => X"d4022800",
		16#4b1a# => X"04000180",
		16#4b1b# => X"9c21fff4",
		16#4b1c# => X"bc2bffff",
		16#4b1d# => X"0c000007",
		16#4b1e# => X"15000000",
		16#4b1f# => X"9c21000c",
		16#4b20# => X"8521fffc",
		16#4b21# => X"8441fff4",
		16#4b22# => X"44004800",
		16#4b23# => X"85c1fff8",
		16#4b24# => X"84420000",
		16#4b25# => X"bc020000",
		16#4b26# => X"13fffff9",
		16#4b27# => X"15000000",
		16#4b28# => X"d40e1000",
		16#4b29# => X"9c21000c",
		16#4b2a# => X"8521fffc",
		16#4b2b# => X"8441fff4",
		16#4b2c# => X"44004800",
		16#4b2d# => X"85c1fff8",
		16#4b2e# => X"d7e117f4",
		16#4b2f# => X"18400001",
		16#4b30# => X"d7e177f8",
		16#4b31# => X"a8429ad0",
		16#4b32# => X"a9c30000",
		16#4b33# => X"a8640000",
		16#4b34# => X"9c800000",
		16#4b35# => X"d7e14ffc",
		16#4b36# => X"d4022000",
		16#4b37# => X"040001ee",
		16#4b38# => X"9c21fff4",
		16#4b39# => X"bc2bffff",
		16#4b3a# => X"0c000007",
		16#4b3b# => X"15000000",
		16#4b3c# => X"9c21000c",
		16#4b3d# => X"8521fffc",
		16#4b3e# => X"8441fff4",
		16#4b3f# => X"44004800",
		16#4b40# => X"85c1fff8",
		16#4b41# => X"84420000",
		16#4b42# => X"bc020000",
		16#4b43# => X"13fffff9",
		16#4b44# => X"15000000",
		16#4b45# => X"d40e1000",
		16#4b46# => X"9c21000c",
		16#4b47# => X"8521fffc",
		16#4b48# => X"8441fff4",
		16#4b49# => X"44004800",
		16#4b4a# => X"85c1fff8",
		16#4b4b# => X"d7e117f4",
		16#4b4c# => X"18400001",
		16#4b4d# => X"d7e177f8",
		16#4b4e# => X"a8429ad0",
		16#4b4f# => X"a9c30000",
		16#4b50# => X"a8640000",
		16#4b51# => X"a8850000",
		16#4b52# => X"a8a60000",
		16#4b53# => X"9cc00000",
		16#4b54# => X"d7e14ffc",
		16#4b55# => X"d4023000",
		16#4b56# => X"040001f8",
		16#4b57# => X"9c21fff4",
		16#4b58# => X"bc2bffff",
		16#4b59# => X"0c000007",
		16#4b5a# => X"15000000",
		16#4b5b# => X"9c21000c",
		16#4b5c# => X"8521fffc",
		16#4b5d# => X"8441fff4",
		16#4b5e# => X"44004800",
		16#4b5f# => X"85c1fff8",
		16#4b60# => X"84420000",
		16#4b61# => X"bc020000",
		16#4b62# => X"13fffff9",
		16#4b63# => X"15000000",
		16#4b64# => X"d40e1000",
		16#4b65# => X"9c21000c",
		16#4b66# => X"8521fffc",
		16#4b67# => X"8441fff4",
		16#4b68# => X"44004800",
		16#4b69# => X"85c1fff8",
		16#4b6a# => X"d7e117f4",
		16#4b6b# => X"18400001",
		16#4b6c# => X"d7e177f8",
		16#4b6d# => X"a8429ad0",
		16#4b6e# => X"a9c30000",
		16#4b6f# => X"a8640000",
		16#4b70# => X"a8850000",
		16#4b71# => X"a8a60000",
		16#4b72# => X"9cc00000",
		16#4b73# => X"d7e14ffc",
		16#4b74# => X"d4023000",
		16#4b75# => X"040001fb",
		16#4b76# => X"9c21fff4",
		16#4b77# => X"bc2bffff",
		16#4b78# => X"0c000007",
		16#4b79# => X"15000000",
		16#4b7a# => X"9c21000c",
		16#4b7b# => X"8521fffc",
		16#4b7c# => X"8441fff4",
		16#4b7d# => X"44004800",
		16#4b7e# => X"85c1fff8",
		16#4b7f# => X"84420000",
		16#4b80# => X"bc020000",
		16#4b81# => X"13fffff9",
		16#4b82# => X"15000000",
		16#4b83# => X"d40e1000",
		16#4b84# => X"9c21000c",
		16#4b85# => X"8521fffc",
		16#4b86# => X"8441fff4",
		16#4b87# => X"44004800",
		16#4b88# => X"85c1fff8",
		16#4b89# => X"d7e117ec",
		16#4b8a# => X"d7e187f4",
		16#4b8b# => X"d7e197f8",
		16#4b8c# => X"d7e14ffc",
		16#4b8d# => X"d7e177f0",
		16#4b8e# => X"aa030000",
		16#4b8f# => X"9c21ffec",
		16#4b90# => X"aa440000",
		16#4b91# => X"bc030000",
		16#4b92# => X"10000006",
		16#4b93# => X"a8450000",
		16#4b94# => X"84830038",
		16#4b95# => X"bc240000",
		16#4b96# => X"0c00003d",
		16#4b97# => X"15000000",
		16#4b98# => X"98a2000c",
		16#4b99# => X"84820018",
		16#4b9a# => X"a465ffff",
		16#4b9b# => X"d4022008",
		16#4b9c# => X"a4830008",
		16#4b9d# => X"bc040000",
		16#4b9e# => X"1000002b",
		16#4b9f# => X"15000000",
		16#4ba0# => X"84c20010",
		16#4ba1# => X"bc260000",
		16#4ba2# => X"0c000027",
		16#4ba3# => X"15000000",
		16#4ba4# => X"a4632000",
		16#4ba5# => X"bc230000",
		16#4ba6# => X"0c00001d",
		16#4ba7# => X"9c80dfff",
		16#4ba8# => X"84620000",
		16#4ba9# => X"84820014",
		16#4baa# => X"e0c33002",
		16#4bab# => X"e5662000",
		16#4bac# => X"10000038",
		16#4bad# => X"9cc60001",
		16#4bae# => X"84a20008",
		16#4baf# => X"a5d200ff",
		16#4bb0# => X"9ca5ffff",
		16#4bb1# => X"9c830001",
		16#4bb2# => X"d4022808",
		16#4bb3# => X"d8037000",
		16#4bb4# => X"d4022000",
		16#4bb5# => X"84620014",
		16#4bb6# => X"e4033000",
		16#4bb7# => X"10000025",
		16#4bb8# => X"bc2e000a",
		16#4bb9# => X"0c00001e",
		16#4bba# => X"15000000",
		16#4bbb# => X"9c210014",
		16#4bbc# => X"a96e0000",
		16#4bbd# => X"8521fffc",
		16#4bbe# => X"8441ffec",
		16#4bbf# => X"85c1fff0",
		16#4bc0# => X"8601fff4",
		16#4bc1# => X"44004800",
		16#4bc2# => X"8641fff8",
		16#4bc3# => X"84620064",
		16#4bc4# => X"a8a52000",
		16#4bc5# => X"e0632003",
		16#4bc6# => X"dc02280c",
		16#4bc7# => X"03ffffe1",
		16#4bc8# => X"d4021864",
		16#4bc9# => X"a8700000",
		16#4bca# => X"07ffe21c",
		16#4bcb# => X"a8820000",
		16#4bcc# => X"bc2b0000",
		16#4bcd# => X"10000020",
		16#4bce# => X"9dc0ffff",
		16#4bcf# => X"98a2000c",
		16#4bd0# => X"84c20010",
		16#4bd1# => X"03ffffd3",
		16#4bd2# => X"a465ffff",
		16#4bd3# => X"07ffec1b",
		16#4bd4# => X"15000000",
		16#4bd5# => X"03ffffc4",
		16#4bd6# => X"98a2000c",
		16#4bd7# => X"9462000c",
		16#4bd8# => X"a4630001",
		16#4bd9# => X"bc030000",
		16#4bda# => X"13ffffe1",
		16#4bdb# => X"15000000",
		16#4bdc# => X"a8700000",
		16#4bdd# => X"07ffeb03",
		16#4bde# => X"a8820000",
		16#4bdf# => X"bc2b0000",
		16#4be0# => X"0fffffdb",
		16#4be1# => X"15000000",
		16#4be2# => X"03ffffd9",
		16#4be3# => X"9dc0ffff",
		16#4be4# => X"a8700000",
		16#4be5# => X"a8820000",
		16#4be6# => X"07ffeafa",
		16#4be7# => X"9dc0ffff",
		16#4be8# => X"bc2b0000",
		16#4be9# => X"13ffffd2",
		16#4bea# => X"9cc00001",
		16#4beb# => X"03ffffc3",
		16#4bec# => X"84620000",
		16#4bed# => X"9462000c",
		16#4bee# => X"a8630040",
		16#4bef# => X"dc02180c",
		16#4bf0# => X"9c400009",
		16#4bf1# => X"03ffffca",
		16#4bf2# => X"d4101000",
		16#4bf3# => X"a8a40000",
		16#4bf4# => X"a8830000",
		16#4bf5# => X"18600001",
		16#4bf6# => X"d7e14ffc",
		16#4bf7# => X"a86363e0",
		16#4bf8# => X"9c21fffc",
		16#4bf9# => X"84630000",
		16#4bfa# => X"9c210004",
		16#4bfb# => X"8521fffc",
		16#4bfc# => X"03ffff8d",
		16#4bfd# => X"15000000",
		16#4bfe# => X"d7e117e8",
		16#4bff# => X"d7e177ec",
		16#4c00# => X"d7e187f0",
		16#4c01# => X"d7e197f4",
		16#4c02# => X"d7e14ffc",
		16#4c03# => X"d7e1a7f8",
		16#4c04# => X"a8440000",
		16#4c05# => X"9c21ffdc",
		16#4c06# => X"aa030000",
		16#4c07# => X"a9c50000",
		16#4c08# => X"bc240000",
		16#4c09# => X"0c00001a",
		16#4c0a# => X"aa460000",
		16#4c0b# => X"18600001",
		16#4c0c# => X"a8636dd4",
		16#4c0d# => X"07ffefcb",
		16#4c0e# => X"86830000",
		16#4c0f# => X"a8700000",
		16#4c10# => X"a8820000",
		16#4c11# => X"a8ae0000",
		16#4c12# => X"a8cb0000",
		16#4c13# => X"4800a000",
		16#4c14# => X"a8f20000",
		16#4c15# => X"bc2bffff",
		16#4c16# => X"10000005",
		16#4c17# => X"9c400000",
		16#4c18# => X"d4121000",
		16#4c19# => X"9c40008a",
		16#4c1a# => X"d4101000",
		16#4c1b# => X"9c210024",
		16#4c1c# => X"8521fffc",
		16#4c1d# => X"8441ffe8",
		16#4c1e# => X"85c1ffec",
		16#4c1f# => X"8601fff0",
		16#4c20# => X"8641fff4",
		16#4c21# => X"44004800",
		16#4c22# => X"8681fff8",
		16#4c23# => X"18600001",
		16#4c24# => X"a8636dd4",
		16#4c25# => X"07ffefb3",
		16#4c26# => X"85c30000",
		16#4c27# => X"a8700000",
		16#4c28# => X"a8810000",
		16#4c29# => X"a8a20000",
		16#4c2a# => X"a8cb0000",
		16#4c2b# => X"48007000",
		16#4c2c# => X"a8f20000",
		16#4c2d# => X"03ffffe9",
		16#4c2e# => X"bc2bffff",
		16#4c2f# => X"d7e117e4",
		16#4c30# => X"d7e177e8",
		16#4c31# => X"d7e197f0",
		16#4c32# => X"d7e14ffc",
		16#4c33# => X"d7e187ec",
		16#4c34# => X"d7e1a7f4",
		16#4c35# => X"d7e1b7f8",
		16#4c36# => X"a8430000",
		16#4c37# => X"9c21ffd8",
		16#4c38# => X"aa440000",
		16#4c39# => X"bc230000",
		16#4c3a# => X"0c00001f",
		16#4c3b# => X"a9c50000",
		16#4c3c# => X"1a000001",
		16#4c3d# => X"18600001",
		16#4c3e# => X"aa1063e0",
		16#4c3f# => X"a8636dd4",
		16#4c40# => X"86d00000",
		16#4c41# => X"07ffef97",
		16#4c42# => X"86830000",
		16#4c43# => X"a8760000",
		16#4c44# => X"a8820000",
		16#4c45# => X"a8b20000",
		16#4c46# => X"a8cb0000",
		16#4c47# => X"4800a000",
		16#4c48# => X"a8ee0000",
		16#4c49# => X"bc2bffff",
		16#4c4a# => X"10000006",
		16#4c4b# => X"9c600000",
		16#4c4c# => X"84500000",
		16#4c4d# => X"d40e1800",
		16#4c4e# => X"9c60008a",
		16#4c4f# => X"d4021800",
		16#4c50# => X"9c210028",
		16#4c51# => X"8521fffc",
		16#4c52# => X"8441ffe4",
		16#4c53# => X"85c1ffe8",
		16#4c54# => X"8601ffec",
		16#4c55# => X"8641fff0",
		16#4c56# => X"8681fff4",
		16#4c57# => X"44004800",
		16#4c58# => X"86c1fff8",
		16#4c59# => X"1a000001",
		16#4c5a# => X"18600001",
		16#4c5b# => X"aa1063e0",
		16#4c5c# => X"a8636dd4",
		16#4c5d# => X"86900000",
		16#4c5e# => X"07ffef7a",
		16#4c5f# => X"86430000",
		16#4c60# => X"a8740000",
		16#4c61# => X"a8810000",
		16#4c62# => X"a8a20000",
		16#4c63# => X"a8cb0000",
		16#4c64# => X"48009000",
		16#4c65# => X"a8ee0000",
		16#4c66# => X"03ffffe4",
		16#4c67# => X"bc2bffff",
		16#4c68# => X"bc040000",
		16#4c69# => X"10000006",
		16#4c6a# => X"bca500ff",
		16#4c6b# => X"0c000006",
		16#4c6c# => X"15000000",
		16#4c6d# => X"d8042800",
		16#4c6e# => X"9c800001",
		16#4c6f# => X"44004800",
		16#4c70# => X"a9640000",
		16#4c71# => X"9ca0008a",
		16#4c72# => X"9c80ffff",
		16#4c73# => X"03fffffc",
		16#4c74# => X"d4032800",
		16#4c75# => X"d7e187f0",
		16#4c76# => X"aa030000",
		16#4c77# => X"18600001",
		16#4c78# => X"d7e14ffc",
		16#4c79# => X"d7e117e8",
		16#4c7a# => X"d7e177ec",
		16#4c7b# => X"d7e197f4",
		16#4c7c# => X"d7e1a7f8",
		16#4c7d# => X"a8636dd4",
		16#4c7e# => X"9c21ffe8",
		16#4c7f# => X"aa860000",
		16#4c80# => X"a9c40000",
		16#4c81# => X"a8450000",
		16#4c82# => X"07ffef56",
		16#4c83# => X"86430000",
		16#4c84# => X"9c210018",
		16#4c85# => X"a8700000",
		16#4c86# => X"a88e0000",
		16#4c87# => X"a8a20000",
		16#4c88# => X"a8f40000",
		16#4c89# => X"a8cb0000",
		16#4c8a# => X"8521fffc",
		16#4c8b# => X"8441ffe8",
		16#4c8c# => X"85c1ffec",
		16#4c8d# => X"8601fff0",
		16#4c8e# => X"8681fff8",
		16#4c8f# => X"44009000",
		16#4c90# => X"8641fff4",
		16#4c91# => X"15000001",
		16#4c92# => X"00000000",
		16#4c93# => X"15000000",
		16#4c94# => X"18600001",
		16#4c95# => X"9c800009",
		16#4c96# => X"a8639ad0",
		16#4c97# => X"9d60ffff",
		16#4c98# => X"44004800",
		16#4c99# => X"d4032000",
		16#4c9a# => X"e0a01802",
		16#4c9b# => X"e0a51804",
		16#4c9c# => X"bd850000",
		16#4c9d# => X"0c00000c",
		16#4c9e# => X"18a00001",
		16#4c9f# => X"aca30001",
		16#4ca0# => X"e0c02802",
		16#4ca1# => X"e0a62804",
		16#4ca2# => X"bd650000",
		16#4ca3# => X"0c00000f",
		16#4ca4# => X"ac630002",
		16#4ca5# => X"9c602000",
		16#4ca6# => X"9d600000",
		16#4ca7# => X"44004800",
		16#4ca8# => X"d4041804",
		16#4ca9# => X"a8a538fc",
		16#4caa# => X"84a50000",
		16#4cab# => X"e0c02802",
		16#4cac# => X"e0a62804",
		16#4cad# => X"bd850000",
		16#4cae# => X"0ffffff2",
		16#4caf# => X"aca30001",
		16#4cb0# => X"03fffff6",
		16#4cb1# => X"9c602000",
		16#4cb2# => X"e0a01802",
		16#4cb3# => X"e0651804",
		16#4cb4# => X"bd830000",
		16#4cb5# => X"0ffffff1",
		16#4cb6# => X"9c602000",
		16#4cb7# => X"18600001",
		16#4cb8# => X"9c800009",
		16#4cb9# => X"a8639ad0",
		16#4cba# => X"9d60ffff",
		16#4cbb# => X"44004800",
		16#4cbc# => X"d4032000",
		16#4cbd# => X"19000001",
		16#4cbe# => X"9c800000",
		16#4cbf# => X"a90863e0",
		16#4cc0# => X"d7e14ffc",
		16#4cc1# => X"84a80000",
		16#4cc2# => X"d7e117f8",
		16#4cc3# => X"9ce50014",
		16#4cc4# => X"9da502ec",
		16#4cc5# => X"d8072018",
		16#4cc6# => X"9d850354",
		16#4cc7# => X"9d6503bc",
		16#4cc8# => X"84680000",
		16#4cc9# => X"d4056804",
		16#4cca# => X"d4052000",
		16#4ccb# => X"d4056008",
		16#4ccc# => X"d405580c",
		16#4ccd# => X"d4052010",
		16#4cce# => X"18a00001",
		16#4ccf# => X"9cc3007c",
		16#4cd0# => X"a8a53ea4",
		16#4cd1# => X"d4032030",
		16#4cd2# => X"d4032834",
		16#4cd3# => X"d4032038",
		16#4cd4# => X"d403203c",
		16#4cd5# => X"d4032040",
		16#4cd6# => X"d4032044",
		16#4cd7# => X"d4032048",
		16#4cd8# => X"d403204c",
		16#4cd9# => X"d4032050",
		16#4cda# => X"d4032054",
		16#4cdb# => X"d4032058",
		16#4cdc# => X"d403205c",
		16#4cdd# => X"d8032060",
		16#4cde# => X"d4072000",
		16#4cdf# => X"d4072004",
		16#4ce0# => X"d4072008",
		16#4ce1# => X"d407200c",
		16#4ce2# => X"d4072010",
		16#4ce3# => X"d4072014",
		16#4ce4# => X"d4062000",
		16#4ce5# => X"d4062004",
		16#4ce6# => X"d4062008",
		16#4ce7# => X"d406200c",
		16#4ce8# => X"d4062010",
		16#4ce9# => X"9c400000",
		16#4cea# => X"84a80000",
		16#4ceb# => X"9c600001",
		16#4cec# => X"d40520a0",
		16#4ced# => X"d40510a4",
		16#4cee# => X"d40518a8",
		16#4cef# => X"9c60330e",
		16#4cf0# => X"9c40abcd",
		16#4cf1# => X"dc0518ac",
		16#4cf2# => X"9c601234",
		16#4cf3# => X"dc0510ae",
		16#4cf4# => X"dc0518b0",
		16#4cf5# => X"9c40e66d",
		16#4cf6# => X"9c60deec",
		16#4cf7# => X"dc0510b2",
		16#4cf8# => X"dc0518b4",
		16#4cf9# => X"9c400005",
		16#4cfa# => X"9c60000b",
		16#4cfb# => X"dc0510b6",
		16#4cfc# => X"dc0518b8",
		16#4cfd# => X"d40520bc",
		16#4cfe# => X"d40520c0",
		16#4cff# => X"d40520c4",
		16#4d00# => X"d40520c8",
		16#4d01# => X"d40520cc",
		16#4d02# => X"d40520d0",
		16#4d03# => X"d40520f8",
		16#4d04# => X"d40520fc",
		16#4d05# => X"d4052100",
		16#4d06# => X"d4052104",
		16#4d07# => X"d4052108",
		16#4d08# => X"d405210c",
		16#4d09# => X"d4052110",
		16#4d0a# => X"d4052114",
		16#4d0b# => X"d4052118",
		16#4d0c# => X"d405211c",
		16#4d0d# => X"d80520d4",
		16#4d0e# => X"d80520dc",
		16#4d0f# => X"d40520f4",
		16#4d10# => X"9c21fff8",
		16#4d11# => X"d4062014",
		16#4d12# => X"d4062018",
		16#4d13# => X"d406201c",
		16#4d14# => X"d4062020",
		16#4d15# => X"d4052148",
		16#4d16# => X"d405214c",
		16#4d17# => X"d4052150",
		16#4d18# => X"d4052154",
		16#4d19# => X"d40522d4",
		16#4d1a# => X"d40521d4",
		16#4d1b# => X"d40522dc",
		16#4d1c# => X"d40522e0",
		16#4d1d# => X"d40522e4",
		16#4d1e# => X"d40522e8",
		16#4d1f# => X"9c210008",
		16#4d20# => X"9c6502ec",
		16#4d21# => X"8521fffc",
		16#4d22# => X"9ca00138",
		16#4d23# => X"03fff036",
		16#4d24# => X"8441fff8",
		16#4d25# => X"e0801802",
		16#4d26# => X"d7e14ffc",
		16#4d27# => X"e0841804",
		16#4d28# => X"bd840000",
		16#4d29# => X"0c00000d",
		16#4d2a# => X"9c21fffc",
		16#4d2b# => X"ac830002",
		16#4d2c# => X"e0a02002",
		16#4d2d# => X"e0852004",
		16#4d2e# => X"bd640000",
		16#4d2f# => X"0c000013",
		16#4d30# => X"15000000",
		16#4d31# => X"9c800001",
		16#4d32# => X"9c210004",
		16#4d33# => X"8521fffc",
		16#4d34# => X"44004800",
		16#4d35# => X"a9640000",
		16#4d36# => X"18a00001",
		16#4d37# => X"a8a538fc",
		16#4d38# => X"84a50000",
		16#4d39# => X"e0c02802",
		16#4d3a# => X"e0a62804",
		16#4d3b# => X"bd850000",
		16#4d3c# => X"0fffffef",
		16#4d3d# => X"9c800001",
		16#4d3e# => X"9c210004",
		16#4d3f# => X"8521fffc",
		16#4d40# => X"44004800",
		16#4d41# => X"a9640000",
		16#4d42# => X"ac630001",
		16#4d43# => X"e0801802",
		16#4d44# => X"e0641804",
		16#4d45# => X"bd630000",
		16#4d46# => X"13ffffeb",
		16#4d47# => X"15000000",
		16#4d48# => X"040000fa",
		16#4d49# => X"15000000",
		16#4d4a# => X"9c600009",
		16#4d4b# => X"9c80ffff",
		16#4d4c# => X"03ffffe6",
		16#4d4d# => X"d40b1800",
		16#4d4e# => X"e0801802",
		16#4d4f# => X"e0841804",
		16#4d50# => X"bd840000",
		16#4d51# => X"0c00000a",
		16#4d52# => X"18800001",
		16#4d53# => X"ac830002",
		16#4d54# => X"e0a02002",
		16#4d55# => X"e0852004",
		16#4d56# => X"bd640000",
		16#4d57# => X"0c00000e",
		16#4d58# => X"15000000",
		16#4d59# => X"44004800",
		16#4d5a# => X"9d600000",
		16#4d5b# => X"9d600000",
		16#4d5c# => X"a88438fc",
		16#4d5d# => X"84840000",
		16#4d5e# => X"e0a02002",
		16#4d5f# => X"e0852004",
		16#4d60# => X"e5845800",
		16#4d61# => X"0ffffff2",
		16#4d62# => X"15000000",
		16#4d63# => X"44004800",
		16#4d64# => X"15000000",
		16#4d65# => X"ac630001",
		16#4d66# => X"e0801802",
		16#4d67# => X"e0641804",
		16#4d68# => X"bd630000",
		16#4d69# => X"13fffff0",
		16#4d6a# => X"9c800009",
		16#4d6b# => X"18600001",
		16#4d6c# => X"a8639ad0",
		16#4d6d# => X"9d60ffff",
		16#4d6e# => X"44004800",
		16#4d6f# => X"d4032000",
		16#4d70# => X"d7e177f4",
		16#4d71# => X"d7e187f8",
		16#4d72# => X"d7e14ffc",
		16#4d73# => X"d7e117f0",
		16#4d74# => X"aa040000",
		16#4d75# => X"9c21fff0",
		16#4d76# => X"bc230000",
		16#4d77# => X"1000001f",
		16#4d78# => X"a9c50000",
		16#4d79# => X"18400001",
		16#4d7a# => X"a84238fc",
		16#4d7b# => X"84420000",
		16#4d7c# => X"bc020000",
		16#4d7d# => X"10000012",
		16#4d7e# => X"bda50000",
		16#4d7f# => X"0c000008",
		16#4d80# => X"a8430000",
		16#4d81# => X"0000000f",
		16#4d82# => X"9c210010",
		16#4d83# => X"9c420001",
		16#4d84# => X"e54e1000",
		16#4d85# => X"0c00000a",
		16#4d86# => X"15000000",
		16#4d87# => X"04000073",
		16#4d88# => X"15000000",
		16#4d89# => X"b96b0018",
		16#4d8a# => X"e0701000",
		16#4d8b# => X"b96b0098",
		16#4d8c# => X"bc0b000a",
		16#4d8d# => X"0ffffff6",
		16#4d8e# => X"d8035800",
		16#4d8f# => X"9c210010",
		16#4d90# => X"a9620000",
		16#4d91# => X"8521fffc",
		16#4d92# => X"8441fff0",
		16#4d93# => X"85c1fff4",
		16#4d94# => X"44004800",
		16#4d95# => X"8601fff8",
		16#4d96# => X"18600001",
		16#4d97# => X"9c800009",
		16#4d98# => X"a8639ad0",
		16#4d99# => X"9c40ffff",
		16#4d9a# => X"03fffff5",
		16#4d9b# => X"d4032000",
		16#4d9c# => X"18800001",
		16#4d9d# => X"18a00001",
		16#4d9e# => X"a8846dd8",
		16#4d9f# => X"a8a563d8",
		16#4da0# => X"85640000",
		16#4da1# => X"84a50000",
		16#4da2# => X"e06b1800",
		16#4da3# => X"d7e117fc",
		16#4da4# => X"e0a51802",
		16#4da5# => X"18400001",
		16#4da6# => X"e5a51000",
		16#4da7# => X"0c00000a",
		16#4da8# => X"9c21fffc",
		16#4da9# => X"18600001",
		16#4daa# => X"9c80000c",
		16#4dab# => X"a8639ad0",
		16#4dac# => X"9d60ffff",
		16#4dad# => X"d4032000",
		16#4dae# => X"9c210004",
		16#4daf# => X"44004800",
		16#4db0# => X"8441fffc",
		16#4db1# => X"d4041800",
		16#4db2# => X"9c210004",
		16#4db3# => X"44004800",
		16#4db4# => X"8441fffc",
		16#4db5# => X"d7e117f8",
		16#4db6# => X"18400001",
		16#4db7# => X"9c80ffc7",
		16#4db8# => X"a84238fc",
		16#4db9# => X"d7e14ffc",
		16#4dba# => X"84620000",
		16#4dbb# => X"9c21fff8",
		16#4dbc# => X"9c630002",
		16#4dbd# => X"d8032000",
		16#4dbe# => X"9c800000",
		16#4dbf# => X"84620000",
		16#4dc0# => X"9c630001",
		16#4dc1# => X"d8032000",
		16#4dc2# => X"9c800003",
		16#4dc3# => X"84620000",
		16#4dc4# => X"9c630003",
		16#4dc5# => X"d8032000",
		16#4dc6# => X"18600001",
		16#4dc7# => X"18800001",
		16#4dc8# => X"a86338f8",
		16#4dc9# => X"a8843900",
		16#4dca# => X"84630000",
		16#4dcb# => X"07ffc4f6",
		16#4dcc# => X"84840000",
		16#4dcd# => X"84620000",
		16#4dce# => X"9d6b0008",
		16#4dcf# => X"9c630003",
		16#4dd0# => X"b96b0044",
		16#4dd1# => X"8ca30000",
		16#4dd2# => X"a8a50080",
		16#4dd3# => X"a48b00ff",
		16#4dd4# => X"d8032800",
		16#4dd5# => X"b96b0088",
		16#4dd6# => X"84620000",
		16#4dd7# => X"d8032000",
		16#4dd8# => X"a56b00ff",
		16#4dd9# => X"84620000",
		16#4dda# => X"9c630001",
		16#4ddb# => X"d8035800",
		16#4ddc# => X"84420000",
		16#4ddd# => X"9c420003",
		16#4dde# => X"8c620000",
		16#4ddf# => X"a463007f",
		16#4de0# => X"d8021800",
		16#4de1# => X"9c210008",
		16#4de2# => X"8521fffc",
		16#4de3# => X"44004800",
		16#4de4# => X"8441fff8",
		16#4de5# => X"18a00001",
		16#4de6# => X"b8630018",
		16#4de7# => X"a8a538fc",
		16#4de8# => X"84c50000",
		16#4de9# => X"b8e30098",
		16#4dea# => X"9c860005",
		16#4deb# => X"8c640000",
		16#4dec# => X"a4630020",
		16#4ded# => X"bc030000",
		16#4dee# => X"13fffffd",
		16#4def# => X"a46700ff",
		16#4df0# => X"d8061800",
		16#4df1# => X"84850000",
		16#4df2# => X"9c840005",
		16#4df3# => X"8c640000",
		16#4df4# => X"a4630060",
		16#4df5# => X"bc230060",
		16#4df6# => X"13fffffd",
		16#4df7# => X"15000000",
		16#4df8# => X"44004800",
		16#4df9# => X"15000000",
		16#4dfa# => X"18600001",
		16#4dfb# => X"a86338fc",
		16#4dfc# => X"84a30000",
		16#4dfd# => X"9c850005",
		16#4dfe# => X"8c640000",
		16#4dff# => X"a4630001",
		16#4e00# => X"bc030000",
		16#4e01# => X"13fffffd",
		16#4e02# => X"15000000",
		16#4e03# => X"8d650000",
		16#4e04# => X"b96b0018",
		16#4e05# => X"44004800",
		16#4e06# => X"b96b0098",
		16#4e07# => X"d7e187f4",
		16#4e08# => X"d7e197f8",
		16#4e09# => X"d7e14ffc",
		16#4e0a# => X"d7e117ec",
		16#4e0b# => X"d7e177f0",
		16#4e0c# => X"9c63ffff",
		16#4e0d# => X"9c21ffec",
		16#4e0e# => X"aa440000",
		16#4e0f# => X"bc430001",
		16#4e10# => X"1000001f",
		16#4e11# => X"aa050000",
		16#4e12# => X"bd450000",
		16#4e13# => X"0c000014",
		16#4e14# => X"19c00001",
		16#4e15# => X"9c400000",
		16#4e16# => X"00000007",
		16#4e17# => X"a9ce38fc",
		16#4e18# => X"15000004",
		16#4e19# => X"9c420001",
		16#4e1a# => X"e5501000",
		16#4e1b# => X"0c00000c",
		16#4e1c# => X"15000000",
		16#4e1d# => X"848e0000",
		16#4e1e# => X"e0721000",
		16#4e1f# => X"bc040000",
		16#4e20# => X"13fffff8",
		16#4e21# => X"90630000",
		16#4e22# => X"07ffffc3",
		16#4e23# => X"9c420001",
		16#4e24# => X"e5501000",
		16#4e25# => X"13fffff8",
		16#4e26# => X"15000000",
		16#4e27# => X"9c210014",
		16#4e28# => X"a9700000",
		16#4e29# => X"8521fffc",
		16#4e2a# => X"8441ffec",
		16#4e2b# => X"85c1fff0",
		16#4e2c# => X"8601fff4",
		16#4e2d# => X"44004800",
		16#4e2e# => X"8641fff8",
		16#4e2f# => X"18400001",
		16#4e30# => X"9c600009",
		16#4e31# => X"a8429ad0",
		16#4e32# => X"9e00ffff",
		16#4e33# => X"d4021800",
		16#4e34# => X"9c210014",
		16#4e35# => X"a9700000",
		16#4e36# => X"8521fffc",
		16#4e37# => X"8441ffec",
		16#4e38# => X"85c1fff0",
		16#4e39# => X"8601fff4",
		16#4e3a# => X"44004800",
		16#4e3b# => X"8641fff8",
		16#4e3c# => X"00000000",
		16#4e3d# => X"00800000",
		16#4e3e# => X"05f5e100",
		16#4e3f# => X"00000000",
		16#4e40# => X"0001c200",
		16#4e41# => X"0000000d",
		16#4e42# => X"18600001",
		16#4e43# => X"a86363e0",
		16#4e44# => X"44004800",
		16#4e45# => X"85630000",
		16#4e46# => X"9c21fffc",
		16#4e47# => X"d4014800",
		16#4e48# => X"07ffc479",
		16#4e49# => X"15000000",
		16#4e4a# => X"9d670000",
		16#4e4b# => X"85210000",
		16#4e4c# => X"44004800",
		16#4e4d# => X"9c210004",
		16#4e4e# => X"9c21fff8",
		16#4e4f# => X"d4014800",
		16#4e50# => X"d4017004",
		16#4e51# => X"9dc00000",
		16#4e52# => X"e5830000",
		16#4e53# => X"0c000004",
		16#4e54# => X"15000000",
		16#4e55# => X"9dc00001",
		16#4e56# => X"e0601802",
		16#4e57# => X"e5840000",
		16#4e58# => X"0c000003",
		16#4e59# => X"15000000",
		16#4e5a# => X"e0802002",
		16#4e5b# => X"07ffc466",
		16#4e5c# => X"15000000",
		16#4e5d# => X"bc0e0001",
		16#4e5e# => X"0c000003",
		16#4e5f# => X"9d670000",
		16#4e60# => X"e1605802",
		16#4e61# => X"85210000",
		16#4e62# => X"85c10004",
		16#4e63# => X"44004800",
		16#4e64# => X"9c210008",
		16#4e65# => X"d7e117f8",
		16#4e66# => X"18400001",
		16#4e67# => X"d7e14ffc",
		16#4e68# => X"a84263c8",
		16#4e69# => X"8462fffc",
		16#4e6a# => X"bc03ffff",
		16#4e6b# => X"10000009",
		16#4e6c# => X"9c21fff8",
		16#4e6d# => X"9c42fffc",
		16#4e6e# => X"48001800",
		16#4e6f# => X"9c42fffc",
		16#4e70# => X"84620000",
		16#4e71# => X"bc23ffff",
		16#4e72# => X"13fffffc",
		16#4e73# => X"15000000",
		16#4e74# => X"9c210008",
		16#4e75# => X"8521fffc",
		16#4e76# => X"44004800",
		16#4e77# => X"8441fff8",
		16#4e78# => X"d7e14ffc",
		16#4e79# => X"9c21fffc",
		16#4e7a# => X"9c210004",
		16#4e7b# => X"8521fffc",
		16#4e7c# => X"44004800",
		16#4e7d# => X"15000000",
		16#4e7e# => X"9c21fffc",
		16#4e7f# => X"d4014800",
		16#4e80# => X"07ffb9b9",
		16#4e81# => X"15000000",
		16#4e82# => X"85210000",
		16#4e83# => X"44004800",
		16#4e84# => X"9c210004",
		16#4e85# => X"0a47656e",
		16#4e86# => X"65726174",
		16#4e87# => X"696e6720",
		16#4e88# => X"72616e64",
		16#4e89# => X"6f6d2061",
		16#4e8a# => X"72726179",
		16#4e8b# => X"206f6620",
		16#4e8c# => X"73697a65",
		16#4e8d# => X"2025642e",
		16#4e8e# => X"2e2e0a00",
		16#4e8f# => X"52616e64",
		16#4e90# => X"6f6d2061",
		16#4e91# => X"72726179",
		16#4e92# => X"2067656e",
		16#4e93# => X"65726174",
		16#4e94# => X"696f6e20",
		16#4e95# => X"6661696c",
		16#4e96# => X"65642e00",
		16#4e97# => X"52616e64",
		16#4e98# => X"6f6d2061",
		16#4e99# => X"72726179",
		16#4e9a# => X"2067656e",
		16#4e9b# => X"65726174",
		16#4e9c# => X"65642e00",
		16#4e9d# => X"52756e6e",
		16#4e9e# => X"696e6720",
		16#4e9f# => X"71756963",
		16#4ea0# => X"6b736f72",
		16#4ea1# => X"74207769",
		16#4ea2# => X"74682025",
		16#4ea3# => X"64204350",
		16#4ea4# => X"55287329",
		16#4ea5# => X"2e2e2e0a",
		16#4ea6# => X"0046696e",
		16#4ea7# => X"69736865",
		16#4ea8# => X"6420736f",
		16#4ea9# => X"7274696e",
		16#4eaa# => X"672e2e2e",
		16#4eab# => X"0020436f",
		16#4eac# => X"72726563",
		16#4ead# => X"74206f70",
		16#4eae# => X"65726174",
		16#4eaf# => X"696f6e20",
		16#4eb0# => X"76657269",
		16#4eb1# => X"66696564",
		16#4eb2# => X"2e002043",
		16#4eb3# => X"6f727265",
		16#4eb4# => X"6374206f",
		16#4eb5# => X"70657261",
		16#4eb6# => X"74696f6e",
		16#4eb7# => X"20636f75",
		16#4eb8# => X"6c64206e",
		16#4eb9# => X"6f742062",
		16#4eba# => X"65207665",
		16#4ebb# => X"72696669",
		16#4ebc# => X"65642e00",
		16#4ebd# => X"54696d65",
		16#4ebe# => X"20656c61",
		16#4ebf# => X"70736564",
		16#4ec0# => X"3a202564",
		16#4ec1# => X"206d730a",
		16#4ec2# => X"00286370",
		16#4ec3# => X"75696420",
		16#4ec4# => X"23256429",
		16#4ec5# => X"202d2d2d",
		16#4ec6# => X"2d2d2d2d",
		16#4ec7# => X"2d2d2d2d",
		16#4ec8# => X"2d2d2d2d",
		16#4ec9# => X"2d2d2d2d",
		16#4eca# => X"2d2d2d2d",
		16#4ecb# => X"2d2d2d2d",
		16#4ecc# => X"2d2d2d2d",
		16#4ecd# => X"2d2d2d2d",
		16#4ece# => X"2d2d2d2d",
		16#4ecf# => X"2d2d2d2d",
		16#4ed0# => X"2d2d2d2d",
		16#4ed1# => X"2d2d2d2d",
		16#4ed2# => X"2d2d2d2d",
		16#4ed3# => X"2d2d2d2d",
		16#4ed4# => X"2d2d2d0a",
		16#4ed5# => X"00286370",
		16#4ed6# => X"75696420",
		16#4ed7# => X"23256429",
		16#4ed8# => X"20506572",
		16#4ed9# => X"666f726d",
		16#4eda# => X"616e6365",
		16#4edb# => X"20737461",
		16#4edc# => X"74697374",
		16#4edd# => X"6963730a",
		16#4ede# => X"00286370",
		16#4edf# => X"75696420",
		16#4ee0# => X"23256429",
		16#4ee1# => X"20253773",
		16#4ee2# => X"25313173",
		16#4ee3# => X"25347325",
		16#4ee4# => X"38732538",
		16#4ee5# => X"73253132",
		16#4ee6# => X"73253130",
		16#4ee7# => X"730a0045",
		16#4ee8# => X"76656e74",
		16#4ee9# => X"00436f75",
		16#4eea# => X"6e74006d",
		16#4eeb# => X"696e0061",
		16#4eec# => X"7667006d",
		16#4eed# => X"61780054",
		16#4eee# => X"6f74616c",
		16#4eef# => X"00526174",
		16#4ef0# => X"65002863",
		16#4ef1# => X"70756964",
		16#4ef2# => X"20232564",
		16#4ef3# => X"29202537",
		16#4ef4# => X"73253131",
		16#4ef5# => X"75253475",
		16#4ef6# => X"25382e32",
		16#4ef7# => X"66253875",
		16#4ef8# => X"25313275",
		16#4ef9# => X"2531302e",
		16#4efa# => X"35660a00",
		16#4efb# => X"414c5500",
		16#4efc# => X"53484946",
		16#4efd# => X"54004d55",
		16#4efe# => X"4c004a55",
		16#4eff# => X"4d50004f",
		16#4f00# => X"54484552",
		16#4f01# => X"00286370",
		16#4f02# => X"75696420",
		16#4f03# => X"23256429",
		16#4f04# => X"20253773",
		16#4f05# => X"25313175",
		16#4f06# => X"25347525",
		16#4f07# => X"382e3266",
		16#4f08# => X"25387525",
		16#4f09# => X"3132750a",
		16#4f0a# => X"00414c4c",
		16#4f0b# => X"00435248",
		16#4f0c# => X"49465500",
		16#4f0d# => X"43524d49",
		16#4f0e# => X"46550043",
		16#4f0f# => X"52484c53",
		16#4f10# => X"55004352",
		16#4f11# => X"4d4c5355",
		16#4f12# => X"00435748",
		16#4f13# => X"4c535500",
		16#4f14# => X"43574d4c",
		16#4f15# => X"53550028",
		16#4f16# => X"20676c6f",
		16#4f17# => X"62616c20",
		16#4f18# => X"29202d2d",
		16#4f19# => X"2d2d2d2d",
		16#4f1a# => X"2d2d2d2d",
		16#4f1b# => X"2d2d2d2d",
		16#4f1c# => X"2d2d2d2d",
		16#4f1d# => X"2d2d2d2d",
		16#4f1e# => X"2d2d2d2d",
		16#4f1f# => X"2d2d2d2d",
		16#4f20# => X"2d2d2d2d",
		16#4f21# => X"2d2d2d2d",
		16#4f22# => X"2d2d2d2d",
		16#4f23# => X"2d2d2d2d",
		16#4f24# => X"2d2d2d2d",
		16#4f25# => X"2d2d2d2d",
		16#4f26# => X"2d2d2d2d",
		16#4f27# => X"2d2d2d2d",
		16#4f28# => X"00282067",
		16#4f29# => X"6c6f6261",
		16#4f2a# => X"6c202920",
		16#4f2b# => X"476c6f62",
		16#4f2c# => X"616c2070",
		16#4f2d# => X"6572666f",
		16#4f2e# => X"726d616e",
		16#4f2f# => X"63652073",
		16#4f30# => X"74617469",
		16#4f31# => X"73746963",
		16#4f32# => X"73002820",
		16#4f33# => X"676c6f62",
		16#4f34# => X"616c2029",
		16#4f35# => X"20253773",
		16#4f36# => X"25313173",
		16#4f37# => X"25347325",
		16#4f38# => X"38732538",
		16#4f39# => X"73253132",
		16#4f3a# => X"73253130",
		16#4f3b# => X"730a0028",
		16#4f3c# => X"20676c6f",
		16#4f3d# => X"62616c20",
		16#4f3e# => X"29202537",
		16#4f3f# => X"73253131",
		16#4f40# => X"75253475",
		16#4f41# => X"25382e32",
		16#4f42# => X"66253875",
		16#4f43# => X"25313275",
		16#4f44# => X"2531302e",
		16#4f45# => X"35660a00",
		16#4f46# => X"2820676c",
		16#4f47# => X"6f62616c",
		16#4f48# => X"20292025",
		16#4f49# => X"37732531",
		16#4f4a# => X"31752534",
		16#4f4b# => X"7525382e",
		16#4f4c# => X"32662538",
		16#4f4d# => X"75253132",
		16#4f4e# => X"750a0043",
		16#4f4f# => X"4c460043",
		16#4f50# => X"4c574200",
		16#4f51# => X"28637075",
		16#4f52# => X"69642023",
		16#4f53# => X"25642920",
		16#4f54# => X"25735b25",
		16#4f55# => X"32645d20",
		16#4f56# => X"20202020",
		16#4f57# => X"203a2025",
		16#4f58# => X"640a0069",
		16#4f59# => X"6e736e20",
		16#4f5a# => X"4c4f4144",
		16#4f5b# => X"00696e73",
		16#4f5c# => X"6e205354",
		16#4f5d# => X"4f524500",
		16#4f5e# => X"cf000000",
		16#4f5f# => X"00000000",
		16#4f60# => X"00000000",
		16#4f61# => X"00000000",
		16#4f62# => X"00000000",
		16#4f63# => X"00000000",
		16#4f64# => X"00000000",
		16#4f65# => X"00000000",
		16#4f66# => X"00000000",
		16#4f67# => X"00000000",
		16#4f68# => X"00010202",
		16#4f69# => X"03030303",
		16#4f6a# => X"04040404",
		16#4f6b# => X"04040404",
		16#4f6c# => X"05050505",
		16#4f6d# => X"05050505",
		16#4f6e# => X"05050505",
		16#4f6f# => X"05050505",
		16#4f70# => X"06060606",
		16#4f71# => X"06060606",
		16#4f72# => X"06060606",
		16#4f73# => X"06060606",
		16#4f74# => X"06060606",
		16#4f75# => X"06060606",
		16#4f76# => X"06060606",
		16#4f77# => X"06060606",
		16#4f78# => X"07070707",
		16#4f79# => X"07070707",
		16#4f7a# => X"07070707",
		16#4f7b# => X"07070707",
		16#4f7c# => X"07070707",
		16#4f7d# => X"07070707",
		16#4f7e# => X"07070707",
		16#4f7f# => X"07070707",
		16#4f80# => X"07070707",
		16#4f81# => X"07070707",
		16#4f82# => X"07070707",
		16#4f83# => X"07070707",
		16#4f84# => X"07070707",
		16#4f85# => X"07070707",
		16#4f86# => X"07070707",
		16#4f87# => X"07070707",
		16#4f88# => X"08080808",
		16#4f89# => X"08080808",
		16#4f8a# => X"08080808",
		16#4f8b# => X"08080808",
		16#4f8c# => X"08080808",
		16#4f8d# => X"08080808",
		16#4f8e# => X"08080808",
		16#4f8f# => X"08080808",
		16#4f90# => X"08080808",
		16#4f91# => X"08080808",
		16#4f92# => X"08080808",
		16#4f93# => X"08080808",
		16#4f94# => X"08080808",
		16#4f95# => X"08080808",
		16#4f96# => X"08080808",
		16#4f97# => X"08080808",
		16#4f98# => X"08080808",
		16#4f99# => X"08080808",
		16#4f9a# => X"08080808",
		16#4f9b# => X"08080808",
		16#4f9c# => X"08080808",
		16#4f9d# => X"08080808",
		16#4f9e# => X"08080808",
		16#4f9f# => X"08080808",
		16#4fa0# => X"08080808",
		16#4fa1# => X"08080808",
		16#4fa2# => X"08080808",
		16#4fa3# => X"08080808",
		16#4fa4# => X"08080808",
		16#4fa5# => X"08080808",
		16#4fa6# => X"08080808",
		16#4fa7# => X"08080808",
		16#4fa8# => X"000163e4",
		16#4fa9# => X"4300494e",
		16#4faa# => X"4600696e",
		16#4fab# => X"66004e41",
		16#4fac# => X"4e006e61",
		16#4fad# => X"6e003031",
		16#4fae# => X"32333435",
		16#4faf# => X"36373839",
		16#4fb0# => X"41424344",
		16#4fb1# => X"45460030",
		16#4fb2# => X"31323334",
		16#4fb3# => X"35363738",
		16#4fb4# => X"39616263",
		16#4fb5# => X"64656600",
		16#4fb6# => X"286e756c",
		16#4fb7# => X"6c290030",
		16#4fb8# => X"00000000",
		16#4fb9# => X"00000000",
		16#4fba# => X"00000000",
		16#4fbb# => X"00009e28",
		16#4fbc# => X"0000989c",
		16#4fbd# => X"0000989c",
		16#4fbe# => X"00009e3c",
		16#4fbf# => X"0000989c",
		16#4fc0# => X"0000989c",
		16#4fc1# => X"0000989c",
		16#4fc2# => X"0000989c",
		16#4fc3# => X"0000989c",
		16#4fc4# => X"0000989c",
		16#4fc5# => X"00009a04",
		16#4fc6# => X"00009e4c",
		16#4fc7# => X"0000989c",
		16#4fc8# => X"00009a2c",
		16#4fc9# => X"00009e98",
		16#4fca# => X"0000989c",
		16#4fcb# => X"00009e54",
		16#4fcc# => X"00009e64",
		16#4fcd# => X"00009e64",
		16#4fce# => X"00009e64",
		16#4fcf# => X"00009e64",
		16#4fd0# => X"00009e64",
		16#4fd1# => X"00009e64",
		16#4fd2# => X"00009e64",
		16#4fd3# => X"00009e64",
		16#4fd4# => X"00009e64",
		16#4fd5# => X"0000989c",
		16#4fd6# => X"0000989c",
		16#4fd7# => X"0000989c",
		16#4fd8# => X"0000989c",
		16#4fd9# => X"0000989c",
		16#4fda# => X"0000989c",
		16#4fdb# => X"0000989c",
		16#4fdc# => X"0000989c",
		16#4fdd# => X"0000989c",
		16#4fde# => X"0000989c",
		16#4fdf# => X"00009ba8",
		16#4fe0# => X"00009cd4",
		16#4fe1# => X"0000989c",
		16#4fe2# => X"00009cd4",
		16#4fe3# => X"0000989c",
		16#4fe4# => X"0000989c",
		16#4fe5# => X"0000989c",
		16#4fe6# => X"0000989c",
		16#4fe7# => X"00009db4",
		16#4fe8# => X"0000989c",
		16#4fe9# => X"0000989c",
		16#4fea# => X"0000a150",
		16#4feb# => X"0000989c",
		16#4fec# => X"0000989c",
		16#4fed# => X"0000989c",
		16#4fee# => X"0000989c",
		16#4fef# => X"0000989c",
		16#4ff0# => X"0000a0b8",
		16#4ff1# => X"0000989c",
		16#4ff2# => X"0000989c",
		16#4ff3# => X"0000a100",
		16#4ff4# => X"0000989c",
		16#4ff5# => X"0000989c",
		16#4ff6# => X"0000989c",
		16#4ff7# => X"0000989c",
		16#4ff8# => X"0000989c",
		16#4ff9# => X"0000989c",
		16#4ffa# => X"0000989c",
		16#4ffb# => X"0000989c",
		16#4ffc# => X"0000989c",
		16#4ffd# => X"0000989c",
		16#4ffe# => X"00009dc4",
		16#4fff# => X"00009dfc",
		16#5000# => X"00009cd4",
		16#5001# => X"00009cd4",
		16#5002# => X"00009cd4",
		16#5003# => X"00009ef0",
		16#5004# => X"00009dfc",
		16#5005# => X"0000989c",
		16#5006# => X"0000989c",
		16#5007# => X"00009f00",
		16#5008# => X"0000989c",
		16#5009# => X"00009f10",
		16#500a# => X"0000a198",
		16#500b# => X"00009f44",
		16#500c# => X"0000a0a8",
		16#500d# => X"0000989c",
		16#500e# => X"00009fa4",
		16#500f# => X"0000989c",
		16#5010# => X"0000a1a0",
		16#5011# => X"0000989c",
		16#5012# => X"0000989c",
		16#5013# => X"0000a018",
		16#5014# => X"30303030",
		16#5015# => X"30303030",
		16#5016# => X"30303030",
		16#5017# => X"30303030",
		16#5018# => X"20202020",
		16#5019# => X"20202020",
		16#501a# => X"20202020",
		16#501b# => X"20202020",
		16#501c# => X"496e6669",
		16#501d# => X"6e697479",
		16#501e# => X"004e614e",
		16#501f# => X"00000000",
		16#5020# => X"00000000",
		16#5021# => X"00000000",
		16#5022# => X"3ff80000",
		16#5023# => X"00000000",
		16#5024# => X"3fd287a7",
		16#5025# => X"636f4361",
		16#5026# => X"3fc68a28",
		16#5027# => X"8b60c8b3",
		16#5028# => X"3fd34413",
		16#5029# => X"509f79fb",
		16#502a# => X"3ff00000",
		16#502b# => X"00000000",
		16#502c# => X"40240000",
		16#502d# => X"00000000",
		16#502e# => X"401c0000",
		16#502f# => X"00000000",
		16#5030# => X"40140000",
		16#5031# => X"00000000",
		16#5032# => X"3fe00000",
		16#5033# => X"00000000",
		16#5034# => X"504f5349",
		16#5035# => X"58000000",
		16#5036# => X"00013aab",
		16#5037# => X"00013b54",
		16#5038# => X"00013b54",
		16#5039# => X"00013b54",
		16#503a# => X"00013b54",
		16#503b# => X"00013b54",
		16#503c# => X"00013b54",
		16#503d# => X"00013b54",
		16#503e# => X"00013b54",
		16#503f# => X"00013b54",
		16#5040# => X"7f7f7f7f",
		16#5041# => X"7f7f7f7f",
		16#5042# => X"7f7f7f7f",
		16#5043# => X"7f7f0000",
		16#5044# => X"40240000",
		16#5045# => X"00000000",
		16#5046# => X"3ff00000",
		16#5047# => X"00000000",
		16#5048# => X"40240000",
		16#5049# => X"00000000",
		16#504a# => X"40590000",
		16#504b# => X"00000000",
		16#504c# => X"408f4000",
		16#504d# => X"00000000",
		16#504e# => X"40c38800",
		16#504f# => X"00000000",
		16#5050# => X"40f86a00",
		16#5051# => X"00000000",
		16#5052# => X"412e8480",
		16#5053# => X"00000000",
		16#5054# => X"416312d0",
		16#5055# => X"00000000",
		16#5056# => X"4197d784",
		16#5057# => X"00000000",
		16#5058# => X"41cdcd65",
		16#5059# => X"00000000",
		16#505a# => X"4202a05f",
		16#505b# => X"20000000",
		16#505c# => X"42374876",
		16#505d# => X"e8000000",
		16#505e# => X"426d1a94",
		16#505f# => X"a2000000",
		16#5060# => X"42a2309c",
		16#5061# => X"e5400000",
		16#5062# => X"42d6bcc4",
		16#5063# => X"1e900000",
		16#5064# => X"430c6bf5",
		16#5065# => X"26340000",
		16#5066# => X"4341c379",
		16#5067# => X"37e08000",
		16#5068# => X"43763457",
		16#5069# => X"85d8a000",
		16#506a# => X"43abc16d",
		16#506b# => X"674ec800",
		16#506c# => X"43e158e4",
		16#506d# => X"60913d00",
		16#506e# => X"4415af1d",
		16#506f# => X"78b58c40",
		16#5070# => X"444b1ae4",
		16#5071# => X"d6e2ef50",
		16#5072# => X"4480f0cf",
		16#5073# => X"064dd592",
		16#5074# => X"44b52d02",
		16#5075# => X"c7e14af6",
		16#5076# => X"44ea7843",
		16#5077# => X"79d99db4",
		16#5078# => X"4341c379",
		16#5079# => X"37e08000",
		16#507a# => X"4693b8b5",
		16#507b# => X"b5056e17",
		16#507c# => X"4d384f03",
		16#507d# => X"e93ff9f5",
		16#507e# => X"5a827748",
		16#507f# => X"f9301d32",
		16#5080# => X"75154fdd",
		16#5081# => X"7f73bf3c",
		16#5082# => X"3c9cd2b2",
		16#5083# => X"97d889bc",
		16#5084# => X"3949f623",
		16#5085# => X"d5a8a733",
		16#5086# => X"32a50ffd",
		16#5087# => X"44f4a73d",
		16#5088# => X"255bba08",
		16#5089# => X"cf8c979d",
		16#508a# => X"0ac80628",
		16#508b# => X"64ac6f43",
		16#508c# => X"00000005",
		16#508d# => X"00000019",
		16#508e# => X"0000007d",
		16#508f# => X"00011d64",
		16#5090# => X"000118d4",
		16#5091# => X"000118d4",
		16#5092# => X"00011d5c",
		16#5093# => X"000118d4",
		16#5094# => X"000118d4",
		16#5095# => X"000118d4",
		16#5096# => X"000118d4",
		16#5097# => X"000118d4",
		16#5098# => X"000118d4",
		16#5099# => X"00011b58",
		16#509a# => X"00011b88",
		16#509b# => X"000118d4",
		16#509c# => X"00011b80",
		16#509d# => X"00011b98",
		16#509e# => X"000118d4",
		16#509f# => X"00011b90",
		16#50a0# => X"00011e20",
		16#50a1# => X"00011e20",
		16#50a2# => X"00011e20",
		16#50a3# => X"00011e20",
		16#50a4# => X"00011e20",
		16#50a5# => X"00011e20",
		16#50a6# => X"00011e20",
		16#50a7# => X"00011e20",
		16#50a8# => X"00011e20",
		16#50a9# => X"000118d4",
		16#50aa# => X"000118d4",
		16#50ab# => X"000118d4",
		16#50ac# => X"000118d4",
		16#50ad# => X"000118d4",
		16#50ae# => X"000118d4",
		16#50af# => X"000118d4",
		16#50b0# => X"000118d4",
		16#50b1# => X"000118d4",
		16#50b2# => X"000118d4",
		16#50b3# => X"00011e14",
		16#50b4# => X"000118d4",
		16#50b5# => X"000118d4",
		16#50b6# => X"000118d4",
		16#50b7# => X"000118d4",
		16#50b8# => X"000118d4",
		16#50b9# => X"000118d4",
		16#50ba# => X"000118d4",
		16#50bb# => X"000118d4",
		16#50bc# => X"000118d4",
		16#50bd# => X"000118d4",
		16#50be# => X"00011a20",
		16#50bf# => X"000118d4",
		16#50c0# => X"000118d4",
		16#50c1# => X"000118d4",
		16#50c2# => X"000118d4",
		16#50c3# => X"000118d4",
		16#50c4# => X"00011b1c",
		16#50c5# => X"000118d4",
		16#50c6# => X"000118d4",
		16#50c7# => X"00011e00",
		16#50c8# => X"000118d4",
		16#50c9# => X"000118d4",
		16#50ca# => X"000118d4",
		16#50cb# => X"000118d4",
		16#50cc# => X"000118d4",
		16#50cd# => X"000118d4",
		16#50ce# => X"000118d4",
		16#50cf# => X"000118d4",
		16#50d0# => X"000118d4",
		16#50d1# => X"000118d4",
		16#50d2# => X"00011dd0",
		16#50d3# => X"00011d80",
		16#50d4# => X"000118d4",
		16#50d5# => X"000118d4",
		16#50d6# => X"000118d4",
		16#50d7# => X"00011d78",
		16#50d8# => X"00011d80",
		16#50d9# => X"000118d4",
		16#50da# => X"000118d4",
		16#50db# => X"00011a18",
		16#50dc# => X"000118d4",
		16#50dd# => X"00011bf0",
		16#50de# => X"00011a24",
		16#50df# => X"00011cb0",
		16#50e0# => X"00011a18",
		16#50e1# => X"000118d4",
		16#50e2# => X"00011cf8",
		16#50e3# => X"000118d4",
		16#50e4# => X"00011b20",
		16#50e5# => X"000118d4",
		16#50e6# => X"000118d4",
		16#50e7# => X"00011c28",
		16#50e8# => X"30303030",
		16#50e9# => X"30303030",
		16#50ea# => X"30303030",
		16#50eb# => X"30303030",
		16#50ec# => X"20202020",
		16#50ed# => X"20202020",
		16#50ee# => X"20202020",
		16#50ef# => X"20202020",
		16#50f0# => X"00000000",
		16#50f1# => X"00000000",
		16#50f2# => X"00000000",
		16#50f3# => X"00000000",
		16#50f4# => X"00000000",
		16#50f5# => X"00000000",
		16#50f6# => X"00000000",
		16#50f7# => X"00000000",
		16#50f8# => X"00000000",
		16#50f9# => X"00000000",
		16#50fa# => X"00000000",
		16#50fb# => X"00000000",
		16#50fc# => X"00000000",
		16#50fd# => X"00000000",
		16#50fe# => X"00000000",
		16#50ff# => X"00000000",
		16#5100# => X"00000000",
		16#5101# => X"00000000",
		16#5102# => X"00000000",
		16#5103# => X"00000000",
		16#5104# => X"00000000",
		16#5105# => X"00000000",
		16#5106# => X"00000000",
		16#5107# => X"00000000",
		16#5108# => X"00000000",
		16#5109# => X"00000000",
		16#510a# => X"00000000",
		16#510b# => X"00000000",
		16#510c# => X"00000000",
		16#510d# => X"00000000",
		16#510e# => X"00000000",
		16#510f# => X"00000000",
		16#5110# => X"00000000",
		16#5111# => X"00000000",
		16#5112# => X"00000000",
		16#5113# => X"00000000",
		16#5114# => X"00000000",
		16#5115# => X"00000000",
		16#5116# => X"00000000",
		16#5117# => X"00000000",
		16#5118# => X"00000000",
		16#5119# => X"00000000",
		16#511a# => X"00000000",
		16#511b# => X"00000000",
		16#511c# => X"00000000",
		16#511d# => X"00000000",
		16#511e# => X"00000000",
		16#511f# => X"00000000",
		16#5120# => X"00000000",
		16#5121# => X"00000000",
		16#5122# => X"00000000",
		16#5123# => X"00000000",
		16#5124# => X"00000000",
		16#5125# => X"00000000",
		16#5126# => X"00000000",
		16#5127# => X"00000000",
		16#5128# => X"00000000",
		16#5129# => X"00000000",
		16#512a# => X"00000000",
		16#512b# => X"00000000",
		16#512c# => X"00000000",
		16#512d# => X"00000000",
		16#512e# => X"00000000",
		16#512f# => X"00000000",
		16#5130# => X"00000000",
		16#5131# => X"00000000",
		16#5132# => X"00000000",
		16#5133# => X"00000000",
		16#5134# => X"00000000",
		16#5135# => X"00000000",
		16#5136# => X"00000000",
		16#5137# => X"00000000",
		16#5138# => X"00000000",
		16#5139# => X"00000000",
		16#513a# => X"00000000",
		16#513b# => X"00000000",
		16#513c# => X"00000000",
		16#513d# => X"00000000",
		16#513e# => X"00000000",
		16#513f# => X"00000000",
		16#5140# => X"00000000",
		16#5141# => X"00000000",
		16#5142# => X"00000000",
		16#5143# => X"00000000",
		16#5144# => X"00000000",
		16#5145# => X"00000000",
		16#5146# => X"00000000",
		16#5147# => X"00000000",
		16#5148# => X"00000000",
		16#5149# => X"00000000",
		16#514a# => X"00000000",
		16#514b# => X"00000000",
		16#514c# => X"00000000",
		16#514d# => X"00000000",
		16#514e# => X"00000000",
		16#514f# => X"00000000",
		16#5150# => X"00000000",
		16#5151# => X"00000000",
		16#5152# => X"00000000",
		16#5153# => X"00000000",
		16#5154# => X"00000000",
		16#5155# => X"00000000",
		16#5156# => X"00000000",
		16#5157# => X"00000000",
		16#5158# => X"00000000",
		16#5159# => X"00000000",
		16#515a# => X"00000000",
		16#515b# => X"00000000",
		16#515c# => X"00000000",
		16#515d# => X"00000000",
		16#515e# => X"00000000",
		16#515f# => X"00000000",
		16#5160# => X"00000000",
		16#5161# => X"00000000",
		16#5162# => X"00000000",
		16#5163# => X"00000000",
		16#5164# => X"00000000",
		16#5165# => X"00000000",
		16#5166# => X"00000000",
		16#5167# => X"00000000",
		16#5168# => X"00000000",
		16#5169# => X"00000000",
		16#516a# => X"00000000",
		16#516b# => X"00000000",
		16#516c# => X"00000000",
		16#516d# => X"00000000",
		16#516e# => X"00000000",
		16#516f# => X"00000000",
		16#5170# => X"00000000",
		16#5171# => X"00000000",
		16#5172# => X"00000000",
		16#5173# => X"00000000",
		16#5174# => X"00000000",
		16#5175# => X"00000000",
		16#5176# => X"00000000",
		16#5177# => X"00000000",
		16#5178# => X"00000000",
		16#5179# => X"00000000",
		16#517a# => X"00000000",
		16#517b# => X"00000000",
		16#517c# => X"00000000",
		16#517d# => X"00000000",
		16#517e# => X"00000000",
		16#517f# => X"00000000",
		16#5180# => X"00000000",
		16#5181# => X"00000000",
		16#5182# => X"00000000",
		16#5183# => X"00000000",
		16#5184# => X"00000000",
		16#5185# => X"00000000",
		16#5186# => X"00000000",
		16#5187# => X"00000000",
		16#5188# => X"00000000",
		16#5189# => X"00000000",
		16#518a# => X"00000000",
		16#518b# => X"00000000",
		16#518c# => X"00000000",
		16#518d# => X"00000000",
		16#518e# => X"00000000",
		16#518f# => X"00000000",
		16#5190# => X"00000000",
		16#5191# => X"00000000",
		16#5192# => X"00000000",
		16#5193# => X"00000000",
		16#5194# => X"00000000",
		16#5195# => X"00000000",
		16#5196# => X"00000000",
		16#5197# => X"00000000",
		16#5198# => X"00000000",
		16#5199# => X"00000000",
		16#519a# => X"00000000",
		16#519b# => X"00000000",
		16#519c# => X"00000000",
		16#519d# => X"00000000",
		16#519e# => X"00000000",
		16#519f# => X"00000000",
		16#51a0# => X"00000000",
		16#51a1# => X"00000000",
		16#51a2# => X"00000000",
		16#51a3# => X"00000000",
		16#51a4# => X"00000000",
		16#51a5# => X"00000000",
		16#51a6# => X"00000000",
		16#51a7# => X"00000000",
		16#51a8# => X"00000000",
		16#51a9# => X"00000000",
		16#51aa# => X"00000000",
		16#51ab# => X"00000000",
		16#51ac# => X"00000000",
		16#51ad# => X"00000000",
		16#51ae# => X"00000000",
		16#51af# => X"00000000",
		16#51b0# => X"00000000",
		16#51b1# => X"00000000",
		16#51b2# => X"00000000",
		16#51b3# => X"00000000",
		16#51b4# => X"00000000",
		16#51b5# => X"00000000",
		16#51b6# => X"00000000",
		16#51b7# => X"00000000",
		16#51b8# => X"00000000",
		16#51b9# => X"00000000",
		16#51ba# => X"00000000",
		16#51bb# => X"00000000",
		16#51bc# => X"00000000",
		16#51bd# => X"00000000",
		16#51be# => X"00000000",
		16#51bf# => X"00000000",
		16#51c0# => X"00000000",
		16#51c1# => X"00000000",
		16#51c2# => X"00000000",
		16#51c3# => X"00000000",
		16#51c4# => X"00000000",
		16#51c5# => X"00000000",
		16#51c6# => X"00000000",
		16#51c7# => X"00000000",
		16#51c8# => X"00000000",
		16#51c9# => X"00000000",
		16#51ca# => X"00000000",
		16#51cb# => X"00000000",
		16#51cc# => X"00000000",
		16#51cd# => X"00000000",
		16#51ce# => X"00000000",
		16#51cf# => X"00000000",
		16#51d0# => X"00000000",
		16#51d1# => X"00000000",
		16#51d2# => X"00000000",
		16#51d3# => X"00000000",
		16#51d4# => X"00000000",
		16#51d5# => X"00000000",
		16#51d6# => X"00000000",
		16#51d7# => X"00000000",
		16#51d8# => X"00000000",
		16#51d9# => X"00000000",
		16#51da# => X"00000000",
		16#51db# => X"00000000",
		16#51dc# => X"00000000",
		16#51dd# => X"00000000",
		16#51de# => X"00000000",
		16#51df# => X"00000000",
		16#51e0# => X"00000000",
		16#51e1# => X"00000000",
		16#51e2# => X"00000000",
		16#51e3# => X"00000000",
		16#51e4# => X"00000000",
		16#51e5# => X"00000000",
		16#51e6# => X"00000000",
		16#51e7# => X"00000000",
		16#51e8# => X"00000000",
		16#51e9# => X"00000000",
		16#51ea# => X"00000000",
		16#51eb# => X"00000000",
		16#51ec# => X"00000000",
		16#51ed# => X"00000000",
		16#51ee# => X"00000000",
		16#51ef# => X"00000000",
		16#51f0# => X"00000000",
		16#51f1# => X"00000000",
		16#51f2# => X"00000000",
		16#51f3# => X"00000000",
		16#51f4# => X"00000000",
		16#51f5# => X"00000000",
		16#51f6# => X"00000000",
		16#51f7# => X"00000000",
		16#51f8# => X"00000000",
		16#51f9# => X"00000000",
		16#51fa# => X"00000000",
		16#51fb# => X"00000000",
		16#51fc# => X"00000000",
		16#51fd# => X"00000000",
		16#51fe# => X"00000000",
		16#51ff# => X"00000000",
		16#5200# => X"00000000",
		16#5201# => X"00000000",
		16#5202# => X"00000000",
		16#5203# => X"00000000",
		16#5204# => X"00000000",
		16#5205# => X"00000000",
		16#5206# => X"00000000",
		16#5207# => X"00000000",
		16#5208# => X"00000000",
		16#5209# => X"00000000",
		16#520a# => X"00000000",
		16#520b# => X"00000000",
		16#520c# => X"00000000",
		16#520d# => X"00000000",
		16#520e# => X"00000000",
		16#520f# => X"00000000",
		16#5210# => X"00000000",
		16#5211# => X"00000000",
		16#5212# => X"00000000",
		16#5213# => X"00000000",
		16#5214# => X"00000000",
		16#5215# => X"00000000",
		16#5216# => X"00000000",
		16#5217# => X"00000000",
		16#5218# => X"00000000",
		16#5219# => X"00000000",
		16#521a# => X"00000000",
		16#521b# => X"00000000",
		16#521c# => X"00000000",
		16#521d# => X"00000000",
		16#521e# => X"00000000",
		16#521f# => X"00000000",
		16#5220# => X"00000000",
		16#5221# => X"00000000",
		16#5222# => X"00000000",
		16#5223# => X"00000000",
		16#5224# => X"00000000",
		16#5225# => X"00000000",
		16#5226# => X"00000000",
		16#5227# => X"00000000",
		16#5228# => X"00000000",
		16#5229# => X"00000000",
		16#522a# => X"00000000",
		16#522b# => X"00000000",
		16#522c# => X"00000000",
		16#522d# => X"00000000",
		16#522e# => X"00000000",
		16#522f# => X"00000000",
		16#5230# => X"00000000",
		16#5231# => X"00000000",
		16#5232# => X"00000000",
		16#5233# => X"00000000",
		16#5234# => X"00000000",
		16#5235# => X"00000000",
		16#5236# => X"00000000",
		16#5237# => X"00000000",
		16#5238# => X"00000000",
		16#5239# => X"00000000",
		16#523a# => X"00000000",
		16#523b# => X"00000000",
		16#523c# => X"00000000",
		16#523d# => X"00000000",
		16#523e# => X"00000000",
		16#523f# => X"00000000",
		16#5240# => X"00000000",
		16#5241# => X"00000000",
		16#5242# => X"00000000",
		16#5243# => X"00000000",
		16#5244# => X"00000000",
		16#5245# => X"00000000",
		16#5246# => X"00000000",
		16#5247# => X"00000000",
		16#5248# => X"00000000",
		16#5249# => X"00000000",
		16#524a# => X"00000000",
		16#524b# => X"00000000",
		16#524c# => X"00000000",
		16#524d# => X"00000000",
		16#524e# => X"00000000",
		16#524f# => X"00000000",
		16#5250# => X"00000000",
		16#5251# => X"00000000",
		16#5252# => X"00000000",
		16#5253# => X"00000000",
		16#5254# => X"00000000",
		16#5255# => X"00000000",
		16#5256# => X"00000000",
		16#5257# => X"00000000",
		16#5258# => X"00000000",
		16#5259# => X"00000000",
		16#525a# => X"00000000",
		16#525b# => X"00000000",
		16#525c# => X"00000000",
		16#525d# => X"00000000",
		16#525e# => X"00000000",
		16#525f# => X"00000000",
		16#5260# => X"00000000",
		16#5261# => X"00000000",
		16#5262# => X"00000000",
		16#5263# => X"00000000",
		16#5264# => X"00000000",
		16#5265# => X"00000000",
		16#5266# => X"00000000",
		16#5267# => X"00000000",
		16#5268# => X"00000000",
		16#5269# => X"00000000",
		16#526a# => X"00000000",
		16#526b# => X"00000000",
		16#526c# => X"00000000",
		16#526d# => X"00000000",
		16#526e# => X"00000000",
		16#526f# => X"00000000",
		16#5270# => X"00000000",
		16#5271# => X"00000000",
		16#5272# => X"00000000",
		16#5273# => X"00000000",
		16#5274# => X"00000000",
		16#5275# => X"00000000",
		16#5276# => X"00000000",
		16#5277# => X"00000000",
		16#5278# => X"00000000",
		16#5279# => X"00000000",
		16#527a# => X"00000000",
		16#527b# => X"00000000",
		16#527c# => X"00000000",
		16#527d# => X"00000000",
		16#527e# => X"00000000",
		16#527f# => X"00000000",
		16#5280# => X"00000000",
		16#5281# => X"00000000",
		16#5282# => X"00000000",
		16#5283# => X"00000000",
		16#5284# => X"00000000",
		16#5285# => X"00000000",
		16#5286# => X"00000000",
		16#5287# => X"00000000",
		16#5288# => X"00000000",
		16#5289# => X"00000000",
		16#528a# => X"00000000",
		16#528b# => X"00000000",
		16#528c# => X"00000000",
		16#528d# => X"00000000",
		16#528e# => X"00000000",
		16#528f# => X"00000000",
		16#5290# => X"00000000",
		16#5291# => X"00000000",
		16#5292# => X"00000000",
		16#5293# => X"00000000",
		16#5294# => X"00000000",
		16#5295# => X"00000000",
		16#5296# => X"00000000",
		16#5297# => X"00000000",
		16#5298# => X"00000000",
		16#5299# => X"00000000",
		16#529a# => X"00000000",
		16#529b# => X"00000000",
		16#529c# => X"00000000",
		16#529d# => X"00000000",
		16#529e# => X"00000000",
		16#529f# => X"00000000",
		16#52a0# => X"00000000",
		16#52a1# => X"00000000",
		16#52a2# => X"00000000",
		16#52a3# => X"00000000",
		16#52a4# => X"00000000",
		16#52a5# => X"00000000",
		16#52a6# => X"00000000",
		16#52a7# => X"00000000",
		16#52a8# => X"00000000",
		16#52a9# => X"00000000",
		16#52aa# => X"00000000",
		16#52ab# => X"00000000",
		16#52ac# => X"00000000",
		16#52ad# => X"00000000",
		16#52ae# => X"00000000",
		16#52af# => X"00000000",
		16#52b0# => X"00000000",
		16#52b1# => X"00000000",
		16#52b2# => X"00000000",
		16#52b3# => X"00000000",
		16#52b4# => X"00000000",
		16#52b5# => X"00000000",
		16#52b6# => X"00000000",
		16#52b7# => X"00000000",
		16#52b8# => X"00000000",
		16#52b9# => X"00000000",
		16#52ba# => X"00000000",
		16#52bb# => X"00000000",
		16#52bc# => X"00000000",
		16#52bd# => X"00000000",
		16#52be# => X"00000000",
		16#52bf# => X"00000000",
		16#52c0# => X"00000000",
		16#52c1# => X"00000000",
		16#52c2# => X"00000000",
		16#52c3# => X"00000000",
		16#52c4# => X"00000000",
		16#52c5# => X"00000000",
		16#52c6# => X"00000000",
		16#52c7# => X"00000000",
		16#52c8# => X"00000000",
		16#52c9# => X"00000000",
		16#52ca# => X"00000000",
		16#52cb# => X"00000000",
		16#52cc# => X"00000000",
		16#52cd# => X"00000000",
		16#52ce# => X"00000000",
		16#52cf# => X"00000000",
		16#52d0# => X"00000000",
		16#52d1# => X"00000000",
		16#52d2# => X"00000000",
		16#52d3# => X"00000000",
		16#52d4# => X"00000000",
		16#52d5# => X"00000000",
		16#52d6# => X"00000000",
		16#52d7# => X"00000000",
		16#52d8# => X"00000000",
		16#52d9# => X"00000000",
		16#52da# => X"00000000",
		16#52db# => X"00000000",
		16#52dc# => X"00000000",
		16#52dd# => X"00000000",
		16#52de# => X"00000000",
		16#52df# => X"00000000",
		16#52e0# => X"00000000",
		16#52e1# => X"00000000",
		16#52e2# => X"00000000",
		16#52e3# => X"00000000",
		16#52e4# => X"00000000",
		16#52e5# => X"00000000",
		16#52e6# => X"00000000",
		16#52e7# => X"00000000",
		16#52e8# => X"00000000",
		16#52e9# => X"00000000",
		16#52ea# => X"00000000",
		16#52eb# => X"00000000",
		16#52ec# => X"00000000",
		16#52ed# => X"00000000",
		16#52ee# => X"00000000",
		16#52ef# => X"00000000",
		16#52f0# => X"00000000",
		16#52f1# => X"00000000",
		16#52f2# => X"00000000",
		16#52f3# => X"00000000",
		16#52f4# => X"00000000",
		16#52f5# => X"00000000",
		16#52f6# => X"00000000",
		16#52f7# => X"00000000",
		16#52f8# => X"00000000",
		16#52f9# => X"00000000",
		16#52fa# => X"00000000",
		16#52fb# => X"00000000",
		16#52fc# => X"00000000",
		16#52fd# => X"00000000",
		16#52fe# => X"00000000",
		16#52ff# => X"00000000",
		16#5300# => X"00000000",
		16#5301# => X"00000000",
		16#5302# => X"00000000",
		16#5303# => X"00000000",
		16#5304# => X"00000000",
		16#5305# => X"00000000",
		16#5306# => X"00000000",
		16#5307# => X"00000000",
		16#5308# => X"00000000",
		16#5309# => X"00000000",
		16#530a# => X"00000000",
		16#530b# => X"00000000",
		16#530c# => X"00000000",
		16#530d# => X"00000000",
		16#530e# => X"00000000",
		16#530f# => X"00000000",
		16#5310# => X"00000000",
		16#5311# => X"00000000",
		16#5312# => X"00000000",
		16#5313# => X"00000000",
		16#5314# => X"00000000",
		16#5315# => X"00000000",
		16#5316# => X"00000000",
		16#5317# => X"00000000",
		16#5318# => X"00000000",
		16#5319# => X"00000000",
		16#531a# => X"00000000",
		16#531b# => X"00000000",
		16#531c# => X"00000000",
		16#531d# => X"00000000",
		16#531e# => X"00000000",
		16#531f# => X"00000000",
		16#5320# => X"00000000",
		16#5321# => X"00000000",
		16#5322# => X"00000000",
		16#5323# => X"00000000",
		16#5324# => X"00000000",
		16#5325# => X"00000000",
		16#5326# => X"00000000",
		16#5327# => X"00000000",
		16#5328# => X"00000000",
		16#5329# => X"00000000",
		16#532a# => X"00000000",
		16#532b# => X"00000000",
		16#532c# => X"00000000",
		16#532d# => X"00000000",
		16#532e# => X"00000000",
		16#532f# => X"00000000",
		16#5330# => X"00000000",
		16#5331# => X"00000000",
		16#5332# => X"00000000",
		16#5333# => X"00000000",
		16#5334# => X"00000000",
		16#5335# => X"00000000",
		16#5336# => X"00000000",
		16#5337# => X"00000000",
		16#5338# => X"00000000",
		16#5339# => X"00000000",
		16#533a# => X"00000000",
		16#533b# => X"00000000",
		16#533c# => X"00000000",
		16#533d# => X"00000000",
		16#533e# => X"00000000",
		16#533f# => X"00000000",
		16#5340# => X"00000000",
		16#5341# => X"00000000",
		16#5342# => X"00000000",
		16#5343# => X"00000000",
		16#5344# => X"00000000",
		16#5345# => X"00000000",
		16#5346# => X"00000000",
		16#5347# => X"00000000",
		16#5348# => X"00000000",
		16#5349# => X"00000000",
		16#534a# => X"00000000",
		16#534b# => X"00000000",
		16#534c# => X"00000000",
		16#534d# => X"00000000",
		16#534e# => X"00000000",
		16#534f# => X"00000000",
		16#5350# => X"00000000",
		16#5351# => X"00000000",
		16#5352# => X"00000000",
		16#5353# => X"00000000",
		16#5354# => X"00000000",
		16#5355# => X"00000000",
		16#5356# => X"00000000",
		16#5357# => X"00000000",
		16#5358# => X"00000000",
		16#5359# => X"00000000",
		16#535a# => X"00000000",
		16#535b# => X"00000000",
		16#535c# => X"00000000",
		16#535d# => X"00000000",
		16#535e# => X"00000000",
		16#535f# => X"00000000",
		16#5360# => X"00000000",
		16#5361# => X"00000000",
		16#5362# => X"00000000",
		16#5363# => X"00000000",
		16#5364# => X"00000000",
		16#5365# => X"00000000",
		16#5366# => X"00000000",
		16#5367# => X"00000000",
		16#5368# => X"00000000",
		16#5369# => X"00000000",
		16#536a# => X"00000000",
		16#536b# => X"00000000",
		16#536c# => X"00000000",
		16#536d# => X"00000000",
		16#536e# => X"00000000",
		16#536f# => X"00000000",
		16#5370# => X"00000000",
		16#5371# => X"00000000",
		16#5372# => X"00000000",
		16#5373# => X"00000000",
		16#5374# => X"00000000",
		16#5375# => X"00000000",
		16#5376# => X"00000000",
		16#5377# => X"00000000",
		16#5378# => X"00000000",
		16#5379# => X"00000000",
		16#537a# => X"00000000",
		16#537b# => X"00000000",
		16#537c# => X"00000000",
		16#537d# => X"00000000",
		16#537e# => X"00000000",
		16#537f# => X"00000000",
		16#5380# => X"00000000",
		16#5381# => X"00000000",
		16#5382# => X"00000000",
		16#5383# => X"00000000",
		16#5384# => X"00000000",
		16#5385# => X"00000000",
		16#5386# => X"00000000",
		16#5387# => X"00000000",
		16#5388# => X"00000000",
		16#5389# => X"00000000",
		16#538a# => X"00000000",
		16#538b# => X"00000000",
		16#538c# => X"00000000",
		16#538d# => X"00000000",
		16#538e# => X"00000000",
		16#538f# => X"00000000",
		16#5390# => X"00000000",
		16#5391# => X"00000000",
		16#5392# => X"00000000",
		16#5393# => X"00000000",
		16#5394# => X"00000000",
		16#5395# => X"00000000",
		16#5396# => X"00000000",
		16#5397# => X"00000000",
		16#5398# => X"00000000",
		16#5399# => X"00000000",
		16#539a# => X"00000000",
		16#539b# => X"00000000",
		16#539c# => X"00000000",
		16#539d# => X"00000000",
		16#539e# => X"00000000",
		16#539f# => X"00000000",
		16#53a0# => X"00000000",
		16#53a1# => X"00000000",
		16#53a2# => X"00000000",
		16#53a3# => X"00000000",
		16#53a4# => X"00000000",
		16#53a5# => X"00000000",
		16#53a6# => X"00000000",
		16#53a7# => X"00000000",
		16#53a8# => X"00000000",
		16#53a9# => X"00000000",
		16#53aa# => X"00000000",
		16#53ab# => X"00000000",
		16#53ac# => X"00000000",
		16#53ad# => X"00000000",
		16#53ae# => X"00000000",
		16#53af# => X"00000000",
		16#53b0# => X"00000000",
		16#53b1# => X"00000000",
		16#53b2# => X"00000000",
		16#53b3# => X"00000000",
		16#53b4# => X"00000000",
		16#53b5# => X"00000000",
		16#53b6# => X"00000000",
		16#53b7# => X"00000000",
		16#53b8# => X"00000000",
		16#53b9# => X"00000000",
		16#53ba# => X"00000000",
		16#53bb# => X"00000000",
		16#53bc# => X"00000000",
		16#53bd# => X"00000000",
		16#53be# => X"00000000",
		16#53bf# => X"00000000",
		16#53c0# => X"00000000",
		16#53c1# => X"00000000",
		16#53c2# => X"00000000",
		16#53c3# => X"00000000",
		16#53c4# => X"00000000",
		16#53c5# => X"00000000",
		16#53c6# => X"00000000",
		16#53c7# => X"00000000",
		16#53c8# => X"00000000",
		16#53c9# => X"00000000",
		16#53ca# => X"00000000",
		16#53cb# => X"00000000",
		16#53cc# => X"00000000",
		16#53cd# => X"00000000",
		16#53ce# => X"00000000",
		16#53cf# => X"00000000",
		16#53d0# => X"00000000",
		16#53d1# => X"00000000",
		16#53d2# => X"00000000",
		16#53d3# => X"00000000",
		16#53d4# => X"00000000",
		16#53d5# => X"00000000",
		16#53d6# => X"00000000",
		16#53d7# => X"00000000",
		16#53d8# => X"00000000",
		16#53d9# => X"00000000",
		16#53da# => X"00000000",
		16#53db# => X"00000000",
		16#53dc# => X"00000000",
		16#53dd# => X"00000000",
		16#53de# => X"00000000",
		16#53df# => X"00000000",
		16#53e0# => X"00000000",
		16#53e1# => X"00000000",
		16#53e2# => X"00000000",
		16#53e3# => X"00000000",
		16#53e4# => X"00000000",
		16#53e5# => X"00000000",
		16#53e6# => X"00000000",
		16#53e7# => X"00000000",
		16#53e8# => X"00000000",
		16#53e9# => X"00000000",
		16#53ea# => X"00000000",
		16#53eb# => X"00000000",
		16#53ec# => X"00000000",
		16#53ed# => X"00000000",
		16#53ee# => X"00000000",
		16#53ef# => X"00000000",
		16#53f0# => X"00000000",
		16#53f1# => X"00000000",
		16#53f2# => X"00000000",
		16#53f3# => X"00000000",
		16#53f4# => X"00000000",
		16#53f5# => X"00000000",
		16#53f6# => X"00000000",
		16#53f7# => X"00000000",
		16#53f8# => X"00000000",
		16#53f9# => X"00000000",
		16#53fa# => X"00000000",
		16#53fb# => X"00000000",
		16#53fc# => X"00000000",
		16#53fd# => X"00000000",
		16#53fe# => X"00000000",
		16#53ff# => X"00000000",
		16#5400# => X"00000000",
		16#5401# => X"00000000",
		16#5402# => X"00000000",
		16#5403# => X"00000000",
		16#5404# => X"00000000",
		16#5405# => X"00000000",
		16#5406# => X"00000000",
		16#5407# => X"00000000",
		16#5408# => X"00000000",
		16#5409# => X"00000000",
		16#540a# => X"00000000",
		16#540b# => X"00000000",
		16#540c# => X"00000000",
		16#540d# => X"00000000",
		16#540e# => X"00000000",
		16#540f# => X"00000000",
		16#5410# => X"00000000",
		16#5411# => X"00000000",
		16#5412# => X"00000000",
		16#5413# => X"00000000",
		16#5414# => X"00000000",
		16#5415# => X"00000000",
		16#5416# => X"00000000",
		16#5417# => X"00000000",
		16#5418# => X"00000000",
		16#5419# => X"00000000",
		16#541a# => X"00000000",
		16#541b# => X"00000000",
		16#541c# => X"00000000",
		16#541d# => X"00000000",
		16#541e# => X"00000000",
		16#541f# => X"00000000",
		16#5420# => X"00000000",
		16#5421# => X"00000000",
		16#5422# => X"00000000",
		16#5423# => X"00000000",
		16#5424# => X"00000000",
		16#5425# => X"00000000",
		16#5426# => X"00000000",
		16#5427# => X"00000000",
		16#5428# => X"00000000",
		16#5429# => X"00000000",
		16#542a# => X"00000000",
		16#542b# => X"00000000",
		16#542c# => X"00000000",
		16#542d# => X"00000000",
		16#542e# => X"00000000",
		16#542f# => X"00000000",
		16#5430# => X"00000000",
		16#5431# => X"00000000",
		16#5432# => X"00000000",
		16#5433# => X"00000000",
		16#5434# => X"00000000",
		16#5435# => X"00000000",
		16#5436# => X"00000000",
		16#5437# => X"00000000",
		16#5438# => X"00000000",
		16#5439# => X"00000000",
		16#543a# => X"00000000",
		16#543b# => X"00000000",
		16#543c# => X"00000000",
		16#543d# => X"00000000",
		16#543e# => X"00000000",
		16#543f# => X"00000000",
		16#5440# => X"00000000",
		16#5441# => X"00000000",
		16#5442# => X"00000000",
		16#5443# => X"00000000",
		16#5444# => X"00000000",
		16#5445# => X"00000000",
		16#5446# => X"00000000",
		16#5447# => X"00000000",
		16#5448# => X"00000000",
		16#5449# => X"00000000",
		16#544a# => X"00000000",
		16#544b# => X"00000000",
		16#544c# => X"00000000",
		16#544d# => X"00000000",
		16#544e# => X"00000000",
		16#544f# => X"00000000",
		16#5450# => X"00000000",
		16#5451# => X"00000000",
		16#5452# => X"00000000",
		16#5453# => X"00000000",
		16#5454# => X"00000000",
		16#5455# => X"00000000",
		16#5456# => X"00000000",
		16#5457# => X"00000000",
		16#5458# => X"00000000",
		16#5459# => X"00000000",
		16#545a# => X"00000000",
		16#545b# => X"00000000",
		16#545c# => X"00000000",
		16#545d# => X"00000000",
		16#545e# => X"00000000",
		16#545f# => X"00000000",
		16#5460# => X"00000000",
		16#5461# => X"00000000",
		16#5462# => X"00000000",
		16#5463# => X"00000000",
		16#5464# => X"00000000",
		16#5465# => X"00000000",
		16#5466# => X"00000000",
		16#5467# => X"00000000",
		16#5468# => X"00000000",
		16#5469# => X"00000000",
		16#546a# => X"00000000",
		16#546b# => X"00000000",
		16#546c# => X"00000000",
		16#546d# => X"00000000",
		16#546e# => X"00000000",
		16#546f# => X"00000000",
		16#5470# => X"00000000",
		16#5471# => X"00000000",
		16#5472# => X"00000000",
		16#5473# => X"00000000",
		16#5474# => X"00000000",
		16#5475# => X"00000000",
		16#5476# => X"00000000",
		16#5477# => X"00000000",
		16#5478# => X"00000000",
		16#5479# => X"00000000",
		16#547a# => X"00000000",
		16#547b# => X"00000000",
		16#547c# => X"00000000",
		16#547d# => X"00000000",
		16#547e# => X"00000000",
		16#547f# => X"00000000",
		16#5480# => X"00000000",
		16#5481# => X"00000000",
		16#5482# => X"00000000",
		16#5483# => X"00000000",
		16#5484# => X"00000000",
		16#5485# => X"00000000",
		16#5486# => X"00000000",
		16#5487# => X"00000000",
		16#5488# => X"00000000",
		16#5489# => X"00000000",
		16#548a# => X"00000000",
		16#548b# => X"00000000",
		16#548c# => X"00000000",
		16#548d# => X"00000000",
		16#548e# => X"00000000",
		16#548f# => X"00000000",
		16#5490# => X"00000000",
		16#5491# => X"00000000",
		16#5492# => X"00000000",
		16#5493# => X"00000000",
		16#5494# => X"00000000",
		16#5495# => X"00000000",
		16#5496# => X"00000000",
		16#5497# => X"00000000",
		16#5498# => X"00000000",
		16#5499# => X"00000000",
		16#549a# => X"00000000",
		16#549b# => X"00000000",
		16#549c# => X"00000000",
		16#549d# => X"00000000",
		16#549e# => X"00000000",
		16#549f# => X"00000000",
		16#54a0# => X"00000000",
		16#54a1# => X"00000000",
		16#54a2# => X"00000000",
		16#54a3# => X"00000000",
		16#54a4# => X"00000000",
		16#54a5# => X"00000000",
		16#54a6# => X"00000000",
		16#54a7# => X"00000000",
		16#54a8# => X"00000000",
		16#54a9# => X"00000000",
		16#54aa# => X"00000000",
		16#54ab# => X"00000000",
		16#54ac# => X"00000000",
		16#54ad# => X"00000000",
		16#54ae# => X"00000000",
		16#54af# => X"00000000",
		16#54b0# => X"00000000",
		16#54b1# => X"00000000",
		16#54b2# => X"00000000",
		16#54b3# => X"00000000",
		16#54b4# => X"00000000",
		16#54b5# => X"00000000",
		16#54b6# => X"00000000",
		16#54b7# => X"00000000",
		16#54b8# => X"00000000",
		16#54b9# => X"00000000",
		16#54ba# => X"00000000",
		16#54bb# => X"00000000",
		16#54bc# => X"00000000",
		16#54bd# => X"00000000",
		16#54be# => X"00000000",
		16#54bf# => X"00000000",
		16#54c0# => X"00000000",
		16#54c1# => X"00000000",
		16#54c2# => X"00000000",
		16#54c3# => X"00000000",
		16#54c4# => X"00000000",
		16#54c5# => X"00000000",
		16#54c6# => X"00000000",
		16#54c7# => X"00000000",
		16#54c8# => X"00000000",
		16#54c9# => X"00000000",
		16#54ca# => X"00000000",
		16#54cb# => X"00000000",
		16#54cc# => X"00000000",
		16#54cd# => X"00000000",
		16#54ce# => X"00000000",
		16#54cf# => X"00000000",
		16#54d0# => X"00000000",
		16#54d1# => X"00000000",
		16#54d2# => X"00000000",
		16#54d3# => X"00000000",
		16#54d4# => X"00000000",
		16#54d5# => X"00000000",
		16#54d6# => X"00000000",
		16#54d7# => X"00000000",
		16#54d8# => X"00000000",
		16#54d9# => X"00000000",
		16#54da# => X"00000000",
		16#54db# => X"00000000",
		16#54dc# => X"00000000",
		16#54dd# => X"00000000",
		16#54de# => X"00000000",
		16#54df# => X"00000000",
		16#54e0# => X"00000000",
		16#54e1# => X"00000000",
		16#54e2# => X"00000000",
		16#54e3# => X"00000000",
		16#54e4# => X"00000000",
		16#54e5# => X"00000000",
		16#54e6# => X"00000000",
		16#54e7# => X"00000000",
		16#54e8# => X"00000000",
		16#54e9# => X"00000000",
		16#54ea# => X"00000000",
		16#54eb# => X"00000000",
		16#54ec# => X"00000000",
		16#54ed# => X"00000000",
		16#54ee# => X"00000000",
		16#54ef# => X"00000000",
		16#54f0# => X"00000000",
		16#54f1# => X"00000000",
		16#54f2# => X"00000000",
		16#54f3# => X"00000000",
		16#54f4# => X"00000000",
		16#54f5# => X"00000000",
		16#54f6# => X"00000000",
		16#54f7# => X"00000000",
		16#54f8# => X"00000000",
		16#54f9# => X"00000000",
		16#54fa# => X"00000000",
		16#54fb# => X"00000000",
		16#54fc# => X"00000000",
		16#54fd# => X"00000000",
		16#54fe# => X"00000000",
		16#54ff# => X"00000000",
		16#5500# => X"00000000",
		16#5501# => X"00000000",
		16#5502# => X"00000000",
		16#5503# => X"00000000",
		16#5504# => X"00000000",
		16#5505# => X"00000000",
		16#5506# => X"00000000",
		16#5507# => X"00000000",
		16#5508# => X"00000000",
		16#5509# => X"00000000",
		16#550a# => X"00000000",
		16#550b# => X"00000000",
		16#550c# => X"00000000",
		16#550d# => X"00000000",
		16#550e# => X"00000000",
		16#550f# => X"00000000",
		16#5510# => X"00000000",
		16#5511# => X"00000000",
		16#5512# => X"00000000",
		16#5513# => X"00000000",
		16#5514# => X"00000000",
		16#5515# => X"00000000",
		16#5516# => X"00000000",
		16#5517# => X"00000000",
		16#5518# => X"00000000",
		16#5519# => X"00000000",
		16#551a# => X"00000000",
		16#551b# => X"00000000",
		16#551c# => X"00000000",
		16#551d# => X"00000000",
		16#551e# => X"00000000",
		16#551f# => X"00000000",
		16#5520# => X"00000000",
		16#5521# => X"00000000",
		16#5522# => X"00000000",
		16#5523# => X"00000000",
		16#5524# => X"00000000",
		16#5525# => X"00000000",
		16#5526# => X"00000000",
		16#5527# => X"00000000",
		16#5528# => X"00000000",
		16#5529# => X"00000000",
		16#552a# => X"00000000",
		16#552b# => X"00000000",
		16#552c# => X"00000000",
		16#552d# => X"00000000",
		16#552e# => X"00000000",
		16#552f# => X"00000000",
		16#5530# => X"00000000",
		16#5531# => X"00000000",
		16#5532# => X"00000000",
		16#5533# => X"00000000",
		16#5534# => X"00000000",
		16#5535# => X"00000000",
		16#5536# => X"00000000",
		16#5537# => X"00000000",
		16#5538# => X"00000000",
		16#5539# => X"00000000",
		16#553a# => X"00000000",
		16#553b# => X"00000000",
		16#553c# => X"00000000",
		16#553d# => X"00000000",
		16#553e# => X"00000000",
		16#553f# => X"00000000",
		16#5540# => X"00000000",
		16#5541# => X"00000000",
		16#5542# => X"00000000",
		16#5543# => X"00000000",
		16#5544# => X"00000000",
		16#5545# => X"00000000",
		16#5546# => X"00000000",
		16#5547# => X"00000000",
		16#5548# => X"00000000",
		16#5549# => X"00000000",
		16#554a# => X"00000000",
		16#554b# => X"00000000",
		16#554c# => X"00000000",
		16#554d# => X"00000000",
		16#554e# => X"00000000",
		16#554f# => X"00000000",
		16#5550# => X"00000000",
		16#5551# => X"00000000",
		16#5552# => X"00000000",
		16#5553# => X"00000000",
		16#5554# => X"00000000",
		16#5555# => X"00000000",
		16#5556# => X"00000000",
		16#5557# => X"00000000",
		16#5558# => X"00000000",
		16#5559# => X"00000000",
		16#555a# => X"00000000",
		16#555b# => X"00000000",
		16#555c# => X"00000000",
		16#555d# => X"00000000",
		16#555e# => X"00000000",
		16#555f# => X"00000000",
		16#5560# => X"00000000",
		16#5561# => X"00000000",
		16#5562# => X"00000000",
		16#5563# => X"00000000",
		16#5564# => X"00000000",
		16#5565# => X"00000000",
		16#5566# => X"00000000",
		16#5567# => X"00000000",
		16#5568# => X"00000000",
		16#5569# => X"00000000",
		16#556a# => X"00000000",
		16#556b# => X"00000000",
		16#556c# => X"00000000",
		16#556d# => X"00000000",
		16#556e# => X"00000000",
		16#556f# => X"00000000",
		16#5570# => X"00000000",
		16#5571# => X"00000000",
		16#5572# => X"00000000",
		16#5573# => X"00000000",
		16#5574# => X"00000000",
		16#5575# => X"00000000",
		16#5576# => X"00000000",
		16#5577# => X"00000000",
		16#5578# => X"00000000",
		16#5579# => X"00000000",
		16#557a# => X"00000000",
		16#557b# => X"00000000",
		16#557c# => X"00000000",
		16#557d# => X"00000000",
		16#557e# => X"00000000",
		16#557f# => X"00000000",
		16#5580# => X"00000000",
		16#5581# => X"00000000",
		16#5582# => X"00000000",
		16#5583# => X"00000000",
		16#5584# => X"00000000",
		16#5585# => X"00000000",
		16#5586# => X"00000000",
		16#5587# => X"00000000",
		16#5588# => X"00000000",
		16#5589# => X"00000000",
		16#558a# => X"00000000",
		16#558b# => X"00000000",
		16#558c# => X"00000000",
		16#558d# => X"00000000",
		16#558e# => X"00000000",
		16#558f# => X"00000000",
		16#5590# => X"00000000",
		16#5591# => X"00000000",
		16#5592# => X"00000000",
		16#5593# => X"00000000",
		16#5594# => X"00000000",
		16#5595# => X"00000000",
		16#5596# => X"00000000",
		16#5597# => X"00000000",
		16#5598# => X"00000000",
		16#5599# => X"00000000",
		16#559a# => X"00000000",
		16#559b# => X"00000000",
		16#559c# => X"00000000",
		16#559d# => X"00000000",
		16#559e# => X"00000000",
		16#559f# => X"00000000",
		16#55a0# => X"00000000",
		16#55a1# => X"00000000",
		16#55a2# => X"00000000",
		16#55a3# => X"00000000",
		16#55a4# => X"00000000",
		16#55a5# => X"00000000",
		16#55a6# => X"00000000",
		16#55a7# => X"00000000",
		16#55a8# => X"00000000",
		16#55a9# => X"00000000",
		16#55aa# => X"00000000",
		16#55ab# => X"00000000",
		16#55ac# => X"00000000",
		16#55ad# => X"00000000",
		16#55ae# => X"00000000",
		16#55af# => X"00000000",
		16#55b0# => X"00000000",
		16#55b1# => X"00000000",
		16#55b2# => X"00000000",
		16#55b3# => X"00000000",
		16#55b4# => X"00000000",
		16#55b5# => X"00000000",
		16#55b6# => X"00000000",
		16#55b7# => X"00000000",
		16#55b8# => X"00000000",
		16#55b9# => X"00000000",
		16#55ba# => X"00000000",
		16#55bb# => X"00000000",
		16#55bc# => X"00000000",
		16#55bd# => X"00000000",
		16#55be# => X"00000000",
		16#55bf# => X"00000000",
		16#55c0# => X"00000000",
		16#55c1# => X"00000000",
		16#55c2# => X"00000000",
		16#55c3# => X"00000000",
		16#55c4# => X"00000000",
		16#55c5# => X"00000000",
		16#55c6# => X"00000000",
		16#55c7# => X"00000000",
		16#55c8# => X"00000000",
		16#55c9# => X"00000000",
		16#55ca# => X"00000000",
		16#55cb# => X"00000000",
		16#55cc# => X"00000000",
		16#55cd# => X"00000000",
		16#55ce# => X"00000000",
		16#55cf# => X"00000000",
		16#55d0# => X"00000000",
		16#55d1# => X"00000000",
		16#55d2# => X"00000000",
		16#55d3# => X"00000000",
		16#55d4# => X"00000000",
		16#55d5# => X"00000000",
		16#55d6# => X"00000000",
		16#55d7# => X"00000000",
		16#55d8# => X"00000000",
		16#55d9# => X"00000000",
		16#55da# => X"00000000",
		16#55db# => X"00000000",
		16#55dc# => X"00000000",
		16#55dd# => X"00000000",
		16#55de# => X"00000000",
		16#55df# => X"00000000",
		16#55e0# => X"00000000",
		16#55e1# => X"00000000",
		16#55e2# => X"00000000",
		16#55e3# => X"00000000",
		16#55e4# => X"00000000",
		16#55e5# => X"00000000",
		16#55e6# => X"00000000",
		16#55e7# => X"00000000",
		16#55e8# => X"00000000",
		16#55e9# => X"00000000",
		16#55ea# => X"00000000",
		16#55eb# => X"00000000",
		16#55ec# => X"00000000",
		16#55ed# => X"00000000",
		16#55ee# => X"00000000",
		16#55ef# => X"00000000",
		16#55f0# => X"00000000",
		16#55f1# => X"00000000",
		16#55f2# => X"00000000",
		16#55f3# => X"00000000",
		16#55f4# => X"00000000",
		16#55f5# => X"00000000",
		16#55f6# => X"00000000",
		16#55f7# => X"00000000",
		16#55f8# => X"00000000",
		16#55f9# => X"00000000",
		16#55fa# => X"00000000",
		16#55fb# => X"00000000",
		16#55fc# => X"00000000",
		16#55fd# => X"00000000",
		16#55fe# => X"00000000",
		16#55ff# => X"00000000",
		16#5600# => X"00000000",
		16#5601# => X"00000000",
		16#5602# => X"00000000",
		16#5603# => X"00000000",
		16#5604# => X"00000000",
		16#5605# => X"00000000",
		16#5606# => X"00000000",
		16#5607# => X"00000000",
		16#5608# => X"00000000",
		16#5609# => X"00000000",
		16#560a# => X"00000000",
		16#560b# => X"00000000",
		16#560c# => X"00000000",
		16#560d# => X"00000000",
		16#560e# => X"00000000",
		16#560f# => X"00000000",
		16#5610# => X"00000000",
		16#5611# => X"00000000",
		16#5612# => X"00000000",
		16#5613# => X"00000000",
		16#5614# => X"00000000",
		16#5615# => X"00000000",
		16#5616# => X"00000000",
		16#5617# => X"00000000",
		16#5618# => X"00000000",
		16#5619# => X"00000000",
		16#561a# => X"00000000",
		16#561b# => X"00000000",
		16#561c# => X"00000000",
		16#561d# => X"00000000",
		16#561e# => X"00000000",
		16#561f# => X"00000000",
		16#5620# => X"00000000",
		16#5621# => X"00000000",
		16#5622# => X"00000000",
		16#5623# => X"00000000",
		16#5624# => X"00000000",
		16#5625# => X"00000000",
		16#5626# => X"00000000",
		16#5627# => X"00000000",
		16#5628# => X"00000000",
		16#5629# => X"00000000",
		16#562a# => X"00000000",
		16#562b# => X"00000000",
		16#562c# => X"00000000",
		16#562d# => X"00000000",
		16#562e# => X"00000000",
		16#562f# => X"00000000",
		16#5630# => X"00000000",
		16#5631# => X"00000000",
		16#5632# => X"00000000",
		16#5633# => X"00000000",
		16#5634# => X"00000000",
		16#5635# => X"00000000",
		16#5636# => X"00000000",
		16#5637# => X"00000000",
		16#5638# => X"00000000",
		16#5639# => X"00000000",
		16#563a# => X"00000000",
		16#563b# => X"00000000",
		16#563c# => X"00000000",
		16#563d# => X"00000000",
		16#563e# => X"00000000",
		16#563f# => X"00000000",
		16#5640# => X"00000000",
		16#5641# => X"00000000",
		16#5642# => X"00000000",
		16#5643# => X"00000000",
		16#5644# => X"00000000",
		16#5645# => X"00000000",
		16#5646# => X"00000000",
		16#5647# => X"00000000",
		16#5648# => X"00000000",
		16#5649# => X"00000000",
		16#564a# => X"00000000",
		16#564b# => X"00000000",
		16#564c# => X"00000000",
		16#564d# => X"00000000",
		16#564e# => X"00000000",
		16#564f# => X"00000000",
		16#5650# => X"00000000",
		16#5651# => X"00000000",
		16#5652# => X"00000000",
		16#5653# => X"00000000",
		16#5654# => X"00000000",
		16#5655# => X"00000000",
		16#5656# => X"00000000",
		16#5657# => X"00000000",
		16#5658# => X"00000000",
		16#5659# => X"00000000",
		16#565a# => X"00000000",
		16#565b# => X"00000000",
		16#565c# => X"00000000",
		16#565d# => X"00000000",
		16#565e# => X"00000000",
		16#565f# => X"00000000",
		16#5660# => X"00000000",
		16#5661# => X"00000000",
		16#5662# => X"00000000",
		16#5663# => X"00000000",
		16#5664# => X"00000000",
		16#5665# => X"00000000",
		16#5666# => X"00000000",
		16#5667# => X"00000000",
		16#5668# => X"00000000",
		16#5669# => X"00000000",
		16#566a# => X"00000000",
		16#566b# => X"00000000",
		16#566c# => X"00000000",
		16#566d# => X"00000000",
		16#566e# => X"00000000",
		16#566f# => X"00000000",
		16#5670# => X"00000000",
		16#5671# => X"00000000",
		16#5672# => X"00000000",
		16#5673# => X"00000000",
		16#5674# => X"00000000",
		16#5675# => X"00000000",
		16#5676# => X"00000000",
		16#5677# => X"00000000",
		16#5678# => X"00000000",
		16#5679# => X"00000000",
		16#567a# => X"00000000",
		16#567b# => X"00000000",
		16#567c# => X"00000000",
		16#567d# => X"00000000",
		16#567e# => X"00000000",
		16#567f# => X"00000000",
		16#5680# => X"00000000",
		16#5681# => X"00000000",
		16#5682# => X"00000000",
		16#5683# => X"00000000",
		16#5684# => X"00000000",
		16#5685# => X"00000000",
		16#5686# => X"00000000",
		16#5687# => X"00000000",
		16#5688# => X"00000000",
		16#5689# => X"00000000",
		16#568a# => X"00000000",
		16#568b# => X"00000000",
		16#568c# => X"00000000",
		16#568d# => X"00000000",
		16#568e# => X"00000000",
		16#568f# => X"00000000",
		16#5690# => X"00000000",
		16#5691# => X"00000000",
		16#5692# => X"00000000",
		16#5693# => X"00000000",
		16#5694# => X"00000000",
		16#5695# => X"00000000",
		16#5696# => X"00000000",
		16#5697# => X"00000000",
		16#5698# => X"00000000",
		16#5699# => X"00000000",
		16#569a# => X"00000000",
		16#569b# => X"00000000",
		16#569c# => X"00000000",
		16#569d# => X"00000000",
		16#569e# => X"00000000",
		16#569f# => X"00000000",
		16#56a0# => X"00000000",
		16#56a1# => X"00000000",
		16#56a2# => X"00000000",
		16#56a3# => X"00000000",
		16#56a4# => X"00000000",
		16#56a5# => X"00000000",
		16#56a6# => X"00000000",
		16#56a7# => X"00000000",
		16#56a8# => X"00000000",
		16#56a9# => X"00000000",
		16#56aa# => X"00000000",
		16#56ab# => X"00000000",
		16#56ac# => X"00000000",
		16#56ad# => X"00000000",
		16#56ae# => X"00000000",
		16#56af# => X"00000000",
		16#56b0# => X"00000000",
		16#56b1# => X"00000000",
		16#56b2# => X"00000000",
		16#56b3# => X"00000000",
		16#56b4# => X"00000000",
		16#56b5# => X"00000000",
		16#56b6# => X"00000000",
		16#56b7# => X"00000000",
		16#56b8# => X"00000000",
		16#56b9# => X"00000000",
		16#56ba# => X"00000000",
		16#56bb# => X"00000000",
		16#56bc# => X"00000000",
		16#56bd# => X"00000000",
		16#56be# => X"00000000",
		16#56bf# => X"00000000",
		16#56c0# => X"00000000",
		16#56c1# => X"00000000",
		16#56c2# => X"00000000",
		16#56c3# => X"00000000",
		16#56c4# => X"00000000",
		16#56c5# => X"00000000",
		16#56c6# => X"00000000",
		16#56c7# => X"00000000",
		16#56c8# => X"00000000",
		16#56c9# => X"00000000",
		16#56ca# => X"00000000",
		16#56cb# => X"00000000",
		16#56cc# => X"00000000",
		16#56cd# => X"00000000",
		16#56ce# => X"00000000",
		16#56cf# => X"00000000",
		16#56d0# => X"00000000",
		16#56d1# => X"00000000",
		16#56d2# => X"00000000",
		16#56d3# => X"00000000",
		16#56d4# => X"00000000",
		16#56d5# => X"00000000",
		16#56d6# => X"00000000",
		16#56d7# => X"00000000",
		16#56d8# => X"00000000",
		16#56d9# => X"00000000",
		16#56da# => X"00000000",
		16#56db# => X"00000000",
		16#56dc# => X"00000000",
		16#56dd# => X"00000000",
		16#56de# => X"00000000",
		16#56df# => X"00000000",
		16#56e0# => X"00000000",
		16#56e1# => X"00000000",
		16#56e2# => X"00000000",
		16#56e3# => X"00000000",
		16#56e4# => X"00000000",
		16#56e5# => X"00000000",
		16#56e6# => X"00000000",
		16#56e7# => X"00000000",
		16#56e8# => X"00000000",
		16#56e9# => X"00000000",
		16#56ea# => X"00000000",
		16#56eb# => X"00000000",
		16#56ec# => X"00000000",
		16#56ed# => X"00000000",
		16#56ee# => X"00000000",
		16#56ef# => X"00000000",
		16#56f0# => X"00000000",
		16#56f1# => X"00000000",
		16#56f2# => X"00000000",
		16#56f3# => X"00000000",
		16#56f4# => X"00000000",
		16#56f5# => X"00000000",
		16#56f6# => X"00000000",
		16#56f7# => X"00000000",
		16#56f8# => X"00000000",
		16#56f9# => X"00000000",
		16#56fa# => X"00000000",
		16#56fb# => X"00000000",
		16#56fc# => X"00000000",
		16#56fd# => X"00000000",
		16#56fe# => X"00000000",
		16#56ff# => X"00000000",
		16#5700# => X"00000000",
		16#5701# => X"00000000",
		16#5702# => X"00000000",
		16#5703# => X"00000000",
		16#5704# => X"00000000",
		16#5705# => X"00000000",
		16#5706# => X"00000000",
		16#5707# => X"00000000",
		16#5708# => X"00000000",
		16#5709# => X"00000000",
		16#570a# => X"00000000",
		16#570b# => X"00000000",
		16#570c# => X"00000000",
		16#570d# => X"00000000",
		16#570e# => X"00000000",
		16#570f# => X"00000000",
		16#5710# => X"00000000",
		16#5711# => X"00000000",
		16#5712# => X"00000000",
		16#5713# => X"00000000",
		16#5714# => X"00000000",
		16#5715# => X"00000000",
		16#5716# => X"00000000",
		16#5717# => X"00000000",
		16#5718# => X"00000000",
		16#5719# => X"00000000",
		16#571a# => X"00000000",
		16#571b# => X"00000000",
		16#571c# => X"00000000",
		16#571d# => X"00000000",
		16#571e# => X"00000000",
		16#571f# => X"00000000",
		16#5720# => X"00000000",
		16#5721# => X"00000000",
		16#5722# => X"00000000",
		16#5723# => X"00000000",
		16#5724# => X"00000000",
		16#5725# => X"00000000",
		16#5726# => X"00000000",
		16#5727# => X"00000000",
		16#5728# => X"00000000",
		16#5729# => X"00000000",
		16#572a# => X"00000000",
		16#572b# => X"00000000",
		16#572c# => X"00000000",
		16#572d# => X"00000000",
		16#572e# => X"00000000",
		16#572f# => X"00000000",
		16#5730# => X"00000000",
		16#5731# => X"00000000",
		16#5732# => X"00000000",
		16#5733# => X"00000000",
		16#5734# => X"00000000",
		16#5735# => X"00000000",
		16#5736# => X"00000000",
		16#5737# => X"00000000",
		16#5738# => X"00000000",
		16#5739# => X"00000000",
		16#573a# => X"00000000",
		16#573b# => X"00000000",
		16#573c# => X"00000000",
		16#573d# => X"00000000",
		16#573e# => X"00000000",
		16#573f# => X"00000000",
		16#5740# => X"00000000",
		16#5741# => X"00000000",
		16#5742# => X"00000000",
		16#5743# => X"00000000",
		16#5744# => X"00000000",
		16#5745# => X"00000000",
		16#5746# => X"00000000",
		16#5747# => X"00000000",
		16#5748# => X"00000000",
		16#5749# => X"00000000",
		16#574a# => X"00000000",
		16#574b# => X"00000000",
		16#574c# => X"00000000",
		16#574d# => X"00000000",
		16#574e# => X"00000000",
		16#574f# => X"00000000",
		16#5750# => X"00000000",
		16#5751# => X"00000000",
		16#5752# => X"00000000",
		16#5753# => X"00000000",
		16#5754# => X"00000000",
		16#5755# => X"00000000",
		16#5756# => X"00000000",
		16#5757# => X"00000000",
		16#5758# => X"00000000",
		16#5759# => X"00000000",
		16#575a# => X"00000000",
		16#575b# => X"00000000",
		16#575c# => X"00000000",
		16#575d# => X"00000000",
		16#575e# => X"00000000",
		16#575f# => X"00000000",
		16#5760# => X"00000000",
		16#5761# => X"00000000",
		16#5762# => X"00000000",
		16#5763# => X"00000000",
		16#5764# => X"00000000",
		16#5765# => X"00000000",
		16#5766# => X"00000000",
		16#5767# => X"00000000",
		16#5768# => X"00000000",
		16#5769# => X"00000000",
		16#576a# => X"00000000",
		16#576b# => X"00000000",
		16#576c# => X"00000000",
		16#576d# => X"00000000",
		16#576e# => X"00000000",
		16#576f# => X"00000000",
		16#5770# => X"00000000",
		16#5771# => X"00000000",
		16#5772# => X"00000000",
		16#5773# => X"00000000",
		16#5774# => X"00000000",
		16#5775# => X"00000000",
		16#5776# => X"00000000",
		16#5777# => X"00000000",
		16#5778# => X"00000000",
		16#5779# => X"00000000",
		16#577a# => X"00000000",
		16#577b# => X"00000000",
		16#577c# => X"00000000",
		16#577d# => X"00000000",
		16#577e# => X"00000000",
		16#577f# => X"00000000",
		16#5780# => X"00000000",
		16#5781# => X"00000000",
		16#5782# => X"00000000",
		16#5783# => X"00000000",
		16#5784# => X"00000000",
		16#5785# => X"00000000",
		16#5786# => X"00000000",
		16#5787# => X"00000000",
		16#5788# => X"00000000",
		16#5789# => X"00000000",
		16#578a# => X"00000000",
		16#578b# => X"00000000",
		16#578c# => X"00000000",
		16#578d# => X"00000000",
		16#578e# => X"00000000",
		16#578f# => X"00000000",
		16#5790# => X"00000000",
		16#5791# => X"00000000",
		16#5792# => X"00000000",
		16#5793# => X"00000000",
		16#5794# => X"00000000",
		16#5795# => X"00000000",
		16#5796# => X"00000000",
		16#5797# => X"00000000",
		16#5798# => X"00000000",
		16#5799# => X"00000000",
		16#579a# => X"00000000",
		16#579b# => X"00000000",
		16#579c# => X"00000000",
		16#579d# => X"00000000",
		16#579e# => X"00000000",
		16#579f# => X"00000000",
		16#57a0# => X"00000000",
		16#57a1# => X"00000000",
		16#57a2# => X"00000000",
		16#57a3# => X"00000000",
		16#57a4# => X"00000000",
		16#57a5# => X"00000000",
		16#57a6# => X"00000000",
		16#57a7# => X"00000000",
		16#57a8# => X"00000000",
		16#57a9# => X"00000000",
		16#57aa# => X"00000000",
		16#57ab# => X"00000000",
		16#57ac# => X"00000000",
		16#57ad# => X"00000000",
		16#57ae# => X"00000000",
		16#57af# => X"00000000",
		16#57b0# => X"00000000",
		16#57b1# => X"00000000",
		16#57b2# => X"00000000",
		16#57b3# => X"00000000",
		16#57b4# => X"00000000",
		16#57b5# => X"00000000",
		16#57b6# => X"00000000",
		16#57b7# => X"00000000",
		16#57b8# => X"00000000",
		16#57b9# => X"00000000",
		16#57ba# => X"00000000",
		16#57bb# => X"00000000",
		16#57bc# => X"00000000",
		16#57bd# => X"00000000",
		16#57be# => X"00000000",
		16#57bf# => X"00000000",
		16#57c0# => X"00000000",
		16#57c1# => X"00000000",
		16#57c2# => X"00000000",
		16#57c3# => X"00000000",
		16#57c4# => X"00000000",
		16#57c5# => X"00000000",
		16#57c6# => X"00000000",
		16#57c7# => X"00000000",
		16#57c8# => X"00000000",
		16#57c9# => X"00000000",
		16#57ca# => X"00000000",
		16#57cb# => X"00000000",
		16#57cc# => X"00000000",
		16#57cd# => X"00000000",
		16#57ce# => X"00000000",
		16#57cf# => X"00000000",
		16#57d0# => X"00000000",
		16#57d1# => X"00000000",
		16#57d2# => X"00000000",
		16#57d3# => X"00000000",
		16#57d4# => X"00000000",
		16#57d5# => X"00000000",
		16#57d6# => X"00000000",
		16#57d7# => X"00000000",
		16#57d8# => X"00000000",
		16#57d9# => X"00000000",
		16#57da# => X"00000000",
		16#57db# => X"00000000",
		16#57dc# => X"00000000",
		16#57dd# => X"00000000",
		16#57de# => X"00000000",
		16#57df# => X"00000000",
		16#57e0# => X"00000000",
		16#57e1# => X"00000000",
		16#57e2# => X"00000000",
		16#57e3# => X"00000000",
		16#57e4# => X"00000000",
		16#57e5# => X"00000000",
		16#57e6# => X"00000000",
		16#57e7# => X"00000000",
		16#57e8# => X"00000000",
		16#57e9# => X"00000000",
		16#57ea# => X"00000000",
		16#57eb# => X"00000000",
		16#57ec# => X"00000000",
		16#57ed# => X"00000000",
		16#57ee# => X"00000000",
		16#57ef# => X"00000000",
		16#57f0# => X"00000000",
		16#57f1# => X"00000000",
		16#57f2# => X"00000000",
		16#57f3# => X"00000000",
		16#57f4# => X"00000000",
		16#57f5# => X"00000000",
		16#57f6# => X"00000000",
		16#57f7# => X"00000000",
		16#57f8# => X"00000000",
		16#57f9# => X"00000000",
		16#57fa# => X"00000000",
		16#57fb# => X"00000000",
		16#57fc# => X"00000000",
		16#57fd# => X"00000000",
		16#57fe# => X"00000000",
		16#57ff# => X"00000000",
		16#5800# => X"00000000",
		16#5801# => X"00000000",
		16#5802# => X"00000000",
		16#5803# => X"00000000",
		16#5804# => X"00000000",
		16#5805# => X"00000000",
		16#5806# => X"00000000",
		16#5807# => X"00000000",
		16#5808# => X"00000000",
		16#5809# => X"00000000",
		16#580a# => X"00000000",
		16#580b# => X"00000000",
		16#580c# => X"00000000",
		16#580d# => X"00000000",
		16#580e# => X"00000000",
		16#580f# => X"00000000",
		16#5810# => X"00000000",
		16#5811# => X"00000000",
		16#5812# => X"00000000",
		16#5813# => X"00000000",
		16#5814# => X"00000000",
		16#5815# => X"00000000",
		16#5816# => X"00000000",
		16#5817# => X"00000000",
		16#5818# => X"00000000",
		16#5819# => X"00000000",
		16#581a# => X"00000000",
		16#581b# => X"00000000",
		16#581c# => X"00000000",
		16#581d# => X"00000000",
		16#581e# => X"00000000",
		16#581f# => X"00000000",
		16#5820# => X"00000000",
		16#5821# => X"00000000",
		16#5822# => X"00000000",
		16#5823# => X"00000000",
		16#5824# => X"00000000",
		16#5825# => X"00000000",
		16#5826# => X"00000000",
		16#5827# => X"00000000",
		16#5828# => X"00000000",
		16#5829# => X"00000000",
		16#582a# => X"00000000",
		16#582b# => X"00000000",
		16#582c# => X"00000000",
		16#582d# => X"00000000",
		16#582e# => X"00000000",
		16#582f# => X"00000000",
		16#5830# => X"00000000",
		16#5831# => X"00000000",
		16#5832# => X"00000000",
		16#5833# => X"00000000",
		16#5834# => X"00000000",
		16#5835# => X"00000000",
		16#5836# => X"00000000",
		16#5837# => X"00000000",
		16#5838# => X"00000000",
		16#5839# => X"00000000",
		16#583a# => X"00000000",
		16#583b# => X"00000000",
		16#583c# => X"00000000",
		16#583d# => X"00000000",
		16#583e# => X"00000000",
		16#583f# => X"00000000",
		16#5840# => X"00000000",
		16#5841# => X"00000000",
		16#5842# => X"00000000",
		16#5843# => X"00000000",
		16#5844# => X"00000000",
		16#5845# => X"00000000",
		16#5846# => X"00000000",
		16#5847# => X"00000000",
		16#5848# => X"00000000",
		16#5849# => X"00000000",
		16#584a# => X"00000000",
		16#584b# => X"00000000",
		16#584c# => X"00000000",
		16#584d# => X"00000000",
		16#584e# => X"00000000",
		16#584f# => X"00000000",
		16#5850# => X"00000000",
		16#5851# => X"00000000",
		16#5852# => X"00000000",
		16#5853# => X"00000000",
		16#5854# => X"00000000",
		16#5855# => X"00000000",
		16#5856# => X"00000000",
		16#5857# => X"00000000",
		16#5858# => X"00000000",
		16#5859# => X"00000000",
		16#585a# => X"00000000",
		16#585b# => X"00000000",
		16#585c# => X"00000000",
		16#585d# => X"00000000",
		16#585e# => X"00000000",
		16#585f# => X"00000000",
		16#5860# => X"00000000",
		16#5861# => X"00000000",
		16#5862# => X"00000000",
		16#5863# => X"00000000",
		16#5864# => X"00000000",
		16#5865# => X"00000000",
		16#5866# => X"00000000",
		16#5867# => X"00000000",
		16#5868# => X"00000000",
		16#5869# => X"00000000",
		16#586a# => X"00000000",
		16#586b# => X"00000000",
		16#586c# => X"00000000",
		16#586d# => X"00000000",
		16#586e# => X"00000000",
		16#586f# => X"00000000",
		16#5870# => X"00000000",
		16#5871# => X"00000000",
		16#5872# => X"00000000",
		16#5873# => X"00000000",
		16#5874# => X"00000000",
		16#5875# => X"00000000",
		16#5876# => X"00000000",
		16#5877# => X"00000000",
		16#5878# => X"00000000",
		16#5879# => X"00000000",
		16#587a# => X"00000000",
		16#587b# => X"00000000",
		16#587c# => X"00000000",
		16#587d# => X"00000000",
		16#587e# => X"00000000",
		16#587f# => X"00000000",
		16#5880# => X"00000000",
		16#5881# => X"00000000",
		16#5882# => X"00000000",
		16#5883# => X"00000000",
		16#5884# => X"00000000",
		16#5885# => X"00000000",
		16#5886# => X"00000000",
		16#5887# => X"00000000",
		16#5888# => X"00000000",
		16#5889# => X"00000000",
		16#588a# => X"00000000",
		16#588b# => X"00000000",
		16#588c# => X"00000000",
		16#588d# => X"00000000",
		16#588e# => X"00000000",
		16#588f# => X"00000000",
		16#5890# => X"00000000",
		16#5891# => X"00000000",
		16#5892# => X"00000000",
		16#5893# => X"00000000",
		16#5894# => X"00000000",
		16#5895# => X"00000000",
		16#5896# => X"00000000",
		16#5897# => X"00000000",
		16#5898# => X"00000000",
		16#5899# => X"00000000",
		16#589a# => X"00000000",
		16#589b# => X"00000000",
		16#589c# => X"00000000",
		16#589d# => X"00000000",
		16#589e# => X"00000000",
		16#589f# => X"00000000",
		16#58a0# => X"00000000",
		16#58a1# => X"00000000",
		16#58a2# => X"00000000",
		16#58a3# => X"00000000",
		16#58a4# => X"00000000",
		16#58a5# => X"00000000",
		16#58a6# => X"00000000",
		16#58a7# => X"00000000",
		16#58a8# => X"00000000",
		16#58a9# => X"00000000",
		16#58aa# => X"00000000",
		16#58ab# => X"00000000",
		16#58ac# => X"00000000",
		16#58ad# => X"00000000",
		16#58ae# => X"00000000",
		16#58af# => X"00000000",
		16#58b0# => X"00000000",
		16#58b1# => X"00000000",
		16#58b2# => X"00000000",
		16#58b3# => X"00000000",
		16#58b4# => X"00000000",
		16#58b5# => X"00000000",
		16#58b6# => X"00000000",
		16#58b7# => X"00000000",
		16#58b8# => X"00000000",
		16#58b9# => X"00000000",
		16#58ba# => X"00000000",
		16#58bb# => X"00000000",
		16#58bc# => X"00000000",
		16#58bd# => X"00000000",
		16#58be# => X"00000000",
		16#58bf# => X"00000000",
		16#58c0# => X"00000000",
		16#58c1# => X"00000000",
		16#58c2# => X"00000000",
		16#58c3# => X"00000000",
		16#58c4# => X"00000000",
		16#58c5# => X"00000000",
		16#58c6# => X"00000000",
		16#58c7# => X"00000000",
		16#58c8# => X"00000000",
		16#58c9# => X"00000000",
		16#58ca# => X"00000000",
		16#58cb# => X"00000000",
		16#58cc# => X"00000000",
		16#58cd# => X"00000000",
		16#58ce# => X"00000000",
		16#58cf# => X"00000000",
		16#58d0# => X"00000000",
		16#58d1# => X"00000000",
		16#58d2# => X"00000000",
		16#58d3# => X"00000000",
		16#58d4# => X"00000000",
		16#58d5# => X"00000000",
		16#58d6# => X"00000000",
		16#58d7# => X"00000000",
		16#58d8# => X"00000000",
		16#58d9# => X"00000000",
		16#58da# => X"00000000",
		16#58db# => X"00000000",
		16#58dc# => X"00000000",
		16#58dd# => X"00000000",
		16#58de# => X"00000000",
		16#58df# => X"00000000",
		16#58e0# => X"00000000",
		16#58e1# => X"00000000",
		16#58e2# => X"00000000",
		16#58e3# => X"00000000",
		16#58e4# => X"00000000",
		16#58e5# => X"00000000",
		16#58e6# => X"00000000",
		16#58e7# => X"00000000",
		16#58e8# => X"00000000",
		16#58e9# => X"00000000",
		16#58ea# => X"00000000",
		16#58eb# => X"00000000",
		16#58ec# => X"00000000",
		16#58ed# => X"00000000",
		16#58ee# => X"00000000",
		16#58ef# => X"00000000",
		16#58f0# => X"00000000",
		16#58f1# => X"ffffffff",
		16#58f2# => X"00000000",
		16#58f3# => X"ffffffff",
		16#58f4# => X"00000000",
		16#58f5# => X"00000000",
		16#58f6# => X"00000000",
		16#58f7# => X"00000000",
		16#58f8# => X"000163e4",
		16#58f9# => X"00000000",
		16#58fa# => X"000166d0",
		16#58fb# => X"00016738",
		16#58fc# => X"000167a0",
		16#58fd# => X"00000000",
		16#58fe# => X"00000000",
		16#58ff# => X"00000000",
		16#5900# => X"00000000",
		16#5901# => X"00000000",
		16#5902# => X"00000000",
		16#5903# => X"00000000",
		16#5904# => X"00000000",
		16#5905# => X"00000000",
		16#5906# => X"00013ea4",
		16#5907# => X"00000000",
		16#5908# => X"00000000",
		16#5909# => X"00000000",
		16#590a# => X"00000000",
		16#590b# => X"00000000",
		16#590c# => X"00000000",
		16#590d# => X"00000000",
		16#590e# => X"00000000",
		16#590f# => X"00000000",
		16#5910# => X"00000000",
		16#5911# => X"00000000",
		16#5912# => X"00000000",
		16#5913# => X"00000000",
		16#5914# => X"00000000",
		16#5915# => X"00000000",
		16#5916# => X"00000000",
		16#5917# => X"00000000",
		16#5918# => X"00000000",
		16#5919# => X"00000000",
		16#591a# => X"00000000",
		16#591b# => X"00000000",
		16#591c# => X"00000000",
		16#591d# => X"00000000",
		16#591e# => X"00000000",
		16#591f# => X"00000000",
		16#5920# => X"00000000",
		16#5921# => X"00000000",
		16#5922# => X"00000000",
		16#5923# => X"00000001",
		16#5924# => X"330eabcd",
		16#5925# => X"1234e66d",
		16#5926# => X"deec0005",
		16#5927# => X"000b0000",
		16#5928# => X"00000000",
		16#5929# => X"00000000",
		16#592a# => X"00000000",
		16#592b# => X"00000000",
		16#592c# => X"00000000",
		16#592d# => X"00000000",
		16#592e# => X"00000000",
		16#592f# => X"00000000",
		16#5930# => X"00000000",
		16#5931# => X"00000000",
		16#5932# => X"00000000",
		16#5933# => X"00000000",
		16#5934# => X"00000000",
		16#5935# => X"00000000",
		16#5936# => X"00000000",
		16#5937# => X"00000000",
		16#5938# => X"00000000",
		16#5939# => X"00000000",
		16#593a# => X"00000000",
		16#593b# => X"00000000",
		16#593c# => X"00000000",
		16#593d# => X"00000000",
		16#593e# => X"00000000",
		16#593f# => X"00000000",
		16#5940# => X"00000000",
		16#5941# => X"00000000",
		16#5942# => X"00000000",
		16#5943# => X"00000000",
		16#5944# => X"00000000",
		16#5945# => X"00000000",
		16#5946# => X"00000000",
		16#5947# => X"00000000",
		16#5948# => X"00000000",
		16#5949# => X"00000000",
		16#594a# => X"00000000",
		16#594b# => X"00000000",
		16#594c# => X"00000000",
		16#594d# => X"00000000",
		16#594e# => X"00000000",
		16#594f# => X"00000000",
		16#5950# => X"00000000",
		16#5951# => X"00000000",
		16#5952# => X"00000000",
		16#5953# => X"00000000",
		16#5954# => X"00000000",
		16#5955# => X"00000000",
		16#5956# => X"00000000",
		16#5957# => X"00000000",
		16#5958# => X"00000000",
		16#5959# => X"00000000",
		16#595a# => X"00000000",
		16#595b# => X"00000000",
		16#595c# => X"00000000",
		16#595d# => X"00000000",
		16#595e# => X"00000000",
		16#595f# => X"00000000",
		16#5960# => X"00000000",
		16#5961# => X"00000000",
		16#5962# => X"00000000",
		16#5963# => X"00000000",
		16#5964# => X"00000000",
		16#5965# => X"00000000",
		16#5966# => X"00000000",
		16#5967# => X"00000000",
		16#5968# => X"00000000",
		16#5969# => X"00000000",
		16#596a# => X"00000000",
		16#596b# => X"00000000",
		16#596c# => X"00000000",
		16#596d# => X"00000000",
		16#596e# => X"00000000",
		16#596f# => X"00000000",
		16#5970# => X"00000000",
		16#5971# => X"00000000",
		16#5972# => X"00000000",
		16#5973# => X"00000000",
		16#5974# => X"00000000",
		16#5975# => X"00000000",
		16#5976# => X"00000000",
		16#5977# => X"00000000",
		16#5978# => X"00000000",
		16#5979# => X"00000000",
		16#597a# => X"00000000",
		16#597b# => X"00000000",
		16#597c# => X"00000000",
		16#597d# => X"00000000",
		16#597e# => X"00000000",
		16#597f# => X"00000000",
		16#5980# => X"00000000",
		16#5981# => X"00000000",
		16#5982# => X"00000000",
		16#5983# => X"00000000",
		16#5984# => X"00000000",
		16#5985# => X"00000000",
		16#5986# => X"00000000",
		16#5987# => X"00000000",
		16#5988# => X"00000000",
		16#5989# => X"00000000",
		16#598a# => X"00000000",
		16#598b# => X"00000000",
		16#598c# => X"00000000",
		16#598d# => X"00000000",
		16#598e# => X"00000000",
		16#598f# => X"00000000",
		16#5990# => X"00000000",
		16#5991# => X"00000000",
		16#5992# => X"00000000",
		16#5993# => X"00000000",
		16#5994# => X"00000000",
		16#5995# => X"00000000",
		16#5996# => X"00000000",
		16#5997# => X"00000000",
		16#5998# => X"00000000",
		16#5999# => X"00000000",
		16#599a# => X"00000000",
		16#599b# => X"00000000",
		16#599c# => X"00000000",
		16#599d# => X"00000000",
		16#599e# => X"00000000",
		16#599f# => X"00000000",
		16#59a0# => X"00000000",
		16#59a1# => X"00000000",
		16#59a2# => X"00000000",
		16#59a3# => X"00000000",
		16#59a4# => X"00000000",
		16#59a5# => X"00000000",
		16#59a6# => X"00000000",
		16#59a7# => X"00000000",
		16#59a8# => X"00000000",
		16#59a9# => X"00000000",
		16#59aa# => X"00000000",
		16#59ab# => X"00000000",
		16#59ac# => X"00000000",
		16#59ad# => X"00000000",
		16#59ae# => X"00000000",
		16#59af# => X"00000000",
		16#59b0# => X"00000000",
		16#59b1# => X"00000000",
		16#59b2# => X"00000000",
		16#59b3# => X"00000000",
		16#59b4# => X"00000000",
		16#59b5# => X"00000000",
		16#59b6# => X"00000000",
		16#59b7# => X"00000000",
		16#59b8# => X"00000000",
		16#59b9# => X"00000000",
		16#59ba# => X"00000000",
		16#59bb# => X"00000000",
		16#59bc# => X"00000000",
		16#59bd# => X"00000000",
		16#59be# => X"00000000",
		16#59bf# => X"00000000",
		16#59c0# => X"00000000",
		16#59c1# => X"00000000",
		16#59c2# => X"00000000",
		16#59c3# => X"00000000",
		16#59c4# => X"00000000",
		16#59c5# => X"00000000",
		16#59c6# => X"00000000",
		16#59c7# => X"00000000",
		16#59c8# => X"00000000",
		16#59c9# => X"00000000",
		16#59ca# => X"00000000",
		16#59cb# => X"00000000",
		16#59cc# => X"00000000",
		16#59cd# => X"00000000",
		16#59ce# => X"00000000",
		16#59cf# => X"00000000",
		16#59d0# => X"00000000",
		16#59d1# => X"00000000",
		16#59d2# => X"00000000",
		16#59d3# => X"00000000",
		16#59d4# => X"00000000",
		16#59d5# => X"00000000",
		16#59d6# => X"00000000",
		16#59d7# => X"00000000",
		16#59d8# => X"00000000",
		16#59d9# => X"00000000",
		16#59da# => X"00000000",
		16#59db# => X"00000000",
		16#59dc# => X"00000000",
		16#59dd# => X"00000000",
		16#59de# => X"00000000",
		16#59df# => X"00000000",
		16#59e0# => X"00000000",
		16#59e1# => X"00000000",
		16#59e2# => X"00000000",
		16#59e3# => X"00000000",
		16#59e4# => X"00000000",
		16#59e5# => X"00000000",
		16#59e6# => X"00000000",
		16#59e7# => X"00000000",
		16#59e8# => X"00000000",
		16#59e9# => X"00000000",
		16#59ea# => X"00000000",
		16#59eb# => X"00000000",
		16#59ec# => X"00000000",
		16#59ed# => X"00000000",
		16#59ee# => X"00000000",
		16#59ef# => X"00000000",
		16#59f0# => X"00000000",
		16#59f1# => X"00000000",
		16#59f2# => X"00000000",
		16#59f3# => X"00000000",
		16#59f4# => X"00000000",
		16#59f5# => X"00000000",
		16#59f6# => X"00000000",
		16#59f7# => X"00000000",
		16#59f8# => X"00000000",
		16#59f9# => X"00000000",
		16#59fa# => X"00000000",
		16#59fb# => X"00000000",
		16#59fc# => X"00000000",
		16#59fd# => X"00000000",
		16#59fe# => X"00000000",
		16#59ff# => X"00000000",
		16#5a00# => X"00000000",
		16#5a01# => X"00000000",
		16#5a02# => X"00000000",
		16#5a03# => X"00000000",
		16#5a04# => X"00016808",
		16#5a05# => X"00016808",
		16#5a06# => X"00016810",
		16#5a07# => X"00016810",
		16#5a08# => X"00016818",
		16#5a09# => X"00016818",
		16#5a0a# => X"00016820",
		16#5a0b# => X"00016820",
		16#5a0c# => X"00016828",
		16#5a0d# => X"00016828",
		16#5a0e# => X"00016830",
		16#5a0f# => X"00016830",
		16#5a10# => X"00016838",
		16#5a11# => X"00016838",
		16#5a12# => X"00016840",
		16#5a13# => X"00016840",
		16#5a14# => X"00016848",
		16#5a15# => X"00016848",
		16#5a16# => X"00016850",
		16#5a17# => X"00016850",
		16#5a18# => X"00016858",
		16#5a19# => X"00016858",
		16#5a1a# => X"00016860",
		16#5a1b# => X"00016860",
		16#5a1c# => X"00016868",
		16#5a1d# => X"00016868",
		16#5a1e# => X"00016870",
		16#5a1f# => X"00016870",
		16#5a20# => X"00016878",
		16#5a21# => X"00016878",
		16#5a22# => X"00016880",
		16#5a23# => X"00016880",
		16#5a24# => X"00016888",
		16#5a25# => X"00016888",
		16#5a26# => X"00016890",
		16#5a27# => X"00016890",
		16#5a28# => X"00016898",
		16#5a29# => X"00016898",
		16#5a2a# => X"000168a0",
		16#5a2b# => X"000168a0",
		16#5a2c# => X"000168a8",
		16#5a2d# => X"000168a8",
		16#5a2e# => X"000168b0",
		16#5a2f# => X"000168b0",
		16#5a30# => X"000168b8",
		16#5a31# => X"000168b8",
		16#5a32# => X"000168c0",
		16#5a33# => X"000168c0",
		16#5a34# => X"000168c8",
		16#5a35# => X"000168c8",
		16#5a36# => X"000168d0",
		16#5a37# => X"000168d0",
		16#5a38# => X"000168d8",
		16#5a39# => X"000168d8",
		16#5a3a# => X"000168e0",
		16#5a3b# => X"000168e0",
		16#5a3c# => X"000168e8",
		16#5a3d# => X"000168e8",
		16#5a3e# => X"000168f0",
		16#5a3f# => X"000168f0",
		16#5a40# => X"000168f8",
		16#5a41# => X"000168f8",
		16#5a42# => X"00016900",
		16#5a43# => X"00016900",
		16#5a44# => X"00016908",
		16#5a45# => X"00016908",
		16#5a46# => X"00016910",
		16#5a47# => X"00016910",
		16#5a48# => X"00016918",
		16#5a49# => X"00016918",
		16#5a4a# => X"00016920",
		16#5a4b# => X"00016920",
		16#5a4c# => X"00016928",
		16#5a4d# => X"00016928",
		16#5a4e# => X"00016930",
		16#5a4f# => X"00016930",
		16#5a50# => X"00016938",
		16#5a51# => X"00016938",
		16#5a52# => X"00016940",
		16#5a53# => X"00016940",
		16#5a54# => X"00016948",
		16#5a55# => X"00016948",
		16#5a56# => X"00016950",
		16#5a57# => X"00016950",
		16#5a58# => X"00016958",
		16#5a59# => X"00016958",
		16#5a5a# => X"00016960",
		16#5a5b# => X"00016960",
		16#5a5c# => X"00016968",
		16#5a5d# => X"00016968",
		16#5a5e# => X"00016970",
		16#5a5f# => X"00016970",
		16#5a60# => X"00016978",
		16#5a61# => X"00016978",
		16#5a62# => X"00016980",
		16#5a63# => X"00016980",
		16#5a64# => X"00016988",
		16#5a65# => X"00016988",
		16#5a66# => X"00016990",
		16#5a67# => X"00016990",
		16#5a68# => X"00016998",
		16#5a69# => X"00016998",
		16#5a6a# => X"000169a0",
		16#5a6b# => X"000169a0",
		16#5a6c# => X"000169a8",
		16#5a6d# => X"000169a8",
		16#5a6e# => X"000169b0",
		16#5a6f# => X"000169b0",
		16#5a70# => X"000169b8",
		16#5a71# => X"000169b8",
		16#5a72# => X"000169c0",
		16#5a73# => X"000169c0",
		16#5a74# => X"000169c8",
		16#5a75# => X"000169c8",
		16#5a76# => X"000169d0",
		16#5a77# => X"000169d0",
		16#5a78# => X"000169d8",
		16#5a79# => X"000169d8",
		16#5a7a# => X"000169e0",
		16#5a7b# => X"000169e0",
		16#5a7c# => X"000169e8",
		16#5a7d# => X"000169e8",
		16#5a7e# => X"000169f0",
		16#5a7f# => X"000169f0",
		16#5a80# => X"000169f8",
		16#5a81# => X"000169f8",
		16#5a82# => X"00016a00",
		16#5a83# => X"00016a00",
		16#5a84# => X"00016a08",
		16#5a85# => X"00016a08",
		16#5a86# => X"00016a10",
		16#5a87# => X"00016a10",
		16#5a88# => X"00016a18",
		16#5a89# => X"00016a18",
		16#5a8a# => X"00016a20",
		16#5a8b# => X"00016a20",
		16#5a8c# => X"00016a28",
		16#5a8d# => X"00016a28",
		16#5a8e# => X"00016a30",
		16#5a8f# => X"00016a30",
		16#5a90# => X"00016a38",
		16#5a91# => X"00016a38",
		16#5a92# => X"00016a40",
		16#5a93# => X"00016a40",
		16#5a94# => X"00016a48",
		16#5a95# => X"00016a48",
		16#5a96# => X"00016a50",
		16#5a97# => X"00016a50",
		16#5a98# => X"00016a58",
		16#5a99# => X"00016a58",
		16#5a9a# => X"00016a60",
		16#5a9b# => X"00016a60",
		16#5a9c# => X"00016a68",
		16#5a9d# => X"00016a68",
		16#5a9e# => X"00016a70",
		16#5a9f# => X"00016a70",
		16#5aa0# => X"00016a78",
		16#5aa1# => X"00016a78",
		16#5aa2# => X"00016a80",
		16#5aa3# => X"00016a80",
		16#5aa4# => X"00016a88",
		16#5aa5# => X"00016a88",
		16#5aa6# => X"00016a90",
		16#5aa7# => X"00016a90",
		16#5aa8# => X"00016a98",
		16#5aa9# => X"00016a98",
		16#5aaa# => X"00016aa0",
		16#5aab# => X"00016aa0",
		16#5aac# => X"00016aa8",
		16#5aad# => X"00016aa8",
		16#5aae# => X"00016ab0",
		16#5aaf# => X"00016ab0",
		16#5ab0# => X"00016ab8",
		16#5ab1# => X"00016ab8",
		16#5ab2# => X"00016ac0",
		16#5ab3# => X"00016ac0",
		16#5ab4# => X"00016ac8",
		16#5ab5# => X"00016ac8",
		16#5ab6# => X"00016ad0",
		16#5ab7# => X"00016ad0",
		16#5ab8# => X"00016ad8",
		16#5ab9# => X"00016ad8",
		16#5aba# => X"00016ae0",
		16#5abb# => X"00016ae0",
		16#5abc# => X"00016ae8",
		16#5abd# => X"00016ae8",
		16#5abe# => X"00016af0",
		16#5abf# => X"00016af0",
		16#5ac0# => X"00016af8",
		16#5ac1# => X"00016af8",
		16#5ac2# => X"00016b00",
		16#5ac3# => X"00016b00",
		16#5ac4# => X"00016b08",
		16#5ac5# => X"00016b08",
		16#5ac6# => X"00016b10",
		16#5ac7# => X"00016b10",
		16#5ac8# => X"00016b18",
		16#5ac9# => X"00016b18",
		16#5aca# => X"00016b20",
		16#5acb# => X"00016b20",
		16#5acc# => X"00016b28",
		16#5acd# => X"00016b28",
		16#5ace# => X"00016b30",
		16#5acf# => X"00016b30",
		16#5ad0# => X"00016b38",
		16#5ad1# => X"00016b38",
		16#5ad2# => X"00016b40",
		16#5ad3# => X"00016b40",
		16#5ad4# => X"00016b48",
		16#5ad5# => X"00016b48",
		16#5ad6# => X"00016b50",
		16#5ad7# => X"00016b50",
		16#5ad8# => X"00016b58",
		16#5ad9# => X"00016b58",
		16#5ada# => X"00016b60",
		16#5adb# => X"00016b60",
		16#5adc# => X"00016b68",
		16#5add# => X"00016b68",
		16#5ade# => X"00016b70",
		16#5adf# => X"00016b70",
		16#5ae0# => X"00016b78",
		16#5ae1# => X"00016b78",
		16#5ae2# => X"00016b80",
		16#5ae3# => X"00016b80",
		16#5ae4# => X"00016b88",
		16#5ae5# => X"00016b88",
		16#5ae6# => X"00016b90",
		16#5ae7# => X"00016b90",
		16#5ae8# => X"00016b98",
		16#5ae9# => X"00016b98",
		16#5aea# => X"00016ba0",
		16#5aeb# => X"00016ba0",
		16#5aec# => X"00016ba8",
		16#5aed# => X"00016ba8",
		16#5aee# => X"00016bb0",
		16#5aef# => X"00016bb0",
		16#5af0# => X"00016bb8",
		16#5af1# => X"00016bb8",
		16#5af2# => X"00016bc0",
		16#5af3# => X"00016bc0",
		16#5af4# => X"00016bc8",
		16#5af5# => X"00016bc8",
		16#5af6# => X"00016bd0",
		16#5af7# => X"00016bd0",
		16#5af8# => X"00016bd8",
		16#5af9# => X"00016bd8",
		16#5afa# => X"00016be0",
		16#5afb# => X"00016be0",
		16#5afc# => X"00016be8",
		16#5afd# => X"00016be8",
		16#5afe# => X"00016bf0",
		16#5aff# => X"00016bf0",
		16#5b00# => X"00016bf8",
		16#5b01# => X"00016bf8",
		16#5b02# => X"00016c00",
		16#5b03# => X"00016c00",
		16#5b04# => X"00020000",
		16#5b05# => X"ffffffff",
		16#5b06# => X"ffffffff",
		16#5b07# => X"ffffffff",
		16#5b08# => X"ffffffff",
		16#5b09# => X"ffffffff",
		16#5b0a# => X"ffffffff",
		16#5b0b# => X"ffffffff",
		16#5b0c# => X"ffffffff",
		16#5b0d# => X"ffffffff",
		16#5b0e# => X"ffffffff",
		16#5b0f# => X"ffffffff",
		16#5b10# => X"ffffffff",
		16#5b11# => X"ffffffff",
		16#5b12# => X"ffffffff",
		16#5b13# => X"ffffffff",
		16#5b14# => X"ffffffff",
		16#5b15# => X"ffffffff",
		16#5b16# => X"ffffffff",
		16#5b17# => X"ffffffff",
		16#5b18# => X"ffffffff",
		16#5b19# => X"ffffffff",
		16#5b1a# => X"ffffffff",
		16#5b1b# => X"ffffffff",
		16#5b1c# => X"ffffffff",
		16#5b1d# => X"ffffffff",
		16#5b1e# => X"ffffffff",
		16#5b1f# => X"ffffffff",
		16#5b20# => X"ffffffff",
		16#5b21# => X"ffffffff",
		16#5b22# => X"ffffffff",
		16#5b23# => X"ffffffff",
		16#5b24# => X"ffffffff",
		16#5b25# => X"ffffffff",
		16#5b26# => X"ffffffff",
		16#5b27# => X"ffffffff",
		16#5b28# => X"ffffffff",
		16#5b29# => X"ffffffff",
		16#5b2a# => X"ffffffff",
		16#5b2b# => X"ffffffff",
		16#5b2c# => X"ffffffff",
		16#5b2d# => X"ffffffff",
		16#5b2e# => X"ffffffff",
		16#5b2f# => X"ffffffff",
		16#5b30# => X"ffffffff",
		16#5b31# => X"ffffffff",
		16#5b32# => X"ffffffff",
		16#5b33# => X"ffffffff",
		16#5b34# => X"ffffffff",
		16#5b35# => X"ffffffff",
		16#5b36# => X"ffffffff",
		16#5b37# => X"ffffffff",
		16#5b38# => X"ffffffff",
		16#5b39# => X"ffffffff",
		16#5b3a# => X"ffffffff",
		16#5b3b# => X"ffffffff",
		16#5b3c# => X"ffffffff",
		16#5b3d# => X"ffffffff",
		16#5b3e# => X"ffffffff",
		16#5b3f# => X"ffffffff",
		16#5b40# => X"ffffffff",
		16#5b41# => X"ffffffff",
		16#5b42# => X"ffffffff",
		16#5b43# => X"ffffffff",
		16#5b44# => X"ffffffff",
		16#5b45# => X"ffffffff",
		16#5b46# => X"ffffffff",
		16#5b47# => X"ffffffff",
		16#5b48# => X"ffffffff",
		16#5b49# => X"ffffffff",
		16#5b4a# => X"ffffffff",
		16#5b4b# => X"ffffffff",
		16#5b4c# => X"ffffffff",
		16#5b4d# => X"ffffffff",
		16#5b4e# => X"ffffffff",
		16#5b4f# => X"ffffffff",
		16#5b50# => X"ffffffff",
		16#5b51# => X"ffffffff",
		16#5b52# => X"ffffffff",
		16#5b53# => X"ffffffff",
		16#5b54# => X"ffffffff",
		16#5b55# => X"ffffffff",
		16#5b56# => X"ffffffff",
		16#5b57# => X"ffffffff",
		16#5b58# => X"ffffffff",
		16#5b59# => X"ffffffff",
		16#5b5a# => X"ffffffff",
		16#5b5b# => X"ffffffff",
		16#5b5c# => X"ffffffff",
		16#5b5d# => X"ffffffff",
		16#5b5e# => X"ffffffff",
		16#5b5f# => X"ffffffff",
		16#5b60# => X"ffffffff",
		16#5b61# => X"ffffffff",
		16#5b62# => X"ffffffff",
		16#5b63# => X"00000001",
		16#5b64# => X"00000001",
		16#5b65# => X"41534349",
		16#5b66# => X"49000000",
		16#5b67# => X"00000000",
		16#5b68# => X"00000000",
		16#5b69# => X"00000000",
		16#5b6a# => X"00000000",
		16#5b6b# => X"00000000",
		16#5b6c# => X"00000000",
		16#5b6d# => X"41534349",
		16#5b6e# => X"49000000",
		16#5b6f# => X"00000000",
		16#5b70# => X"00000000",
		16#5b71# => X"00000000",
		16#5b72# => X"00000000",
		16#5b73# => X"00000000",
		16#5b74# => X"00000000",
		16#5b75# => X"000131a0",
		16#5b76# => X"00019ad4",
		16#5b77# => X"00000000",
		others => X"00000000"
	);

end package;