library ieee;
use ieee.std_logic_1164.all;

library paranut;
use paranut.types.all;

package prog_mem is

	constant PROG_SIZE : integer := 112612;

	constant PROG_DATA : mem_type(0 to PROG_SIZE/4-1) := (
		16#0000# => X"00000000",
		16#0001# => X"00000000",
		16#0002# => X"00000000",
		16#0003# => X"00000000",
		16#0004# => X"00000000",
		16#0005# => X"00000000",
		16#0006# => X"00000000",
		16#0007# => X"00000000",
		16#0008# => X"00000000",
		16#0009# => X"00000000",
		16#000a# => X"00000000",
		16#000b# => X"00000000",
		16#000c# => X"00000000",
		16#000d# => X"00000000",
		16#000e# => X"00000000",
		16#000f# => X"00000000",
		16#0010# => X"00000000",
		16#0011# => X"00000000",
		16#0012# => X"00000000",
		16#0013# => X"00000000",
		16#0014# => X"00000000",
		16#0015# => X"00000000",
		16#0016# => X"00000000",
		16#0017# => X"00000000",
		16#0018# => X"00000000",
		16#0019# => X"00000000",
		16#001a# => X"00000000",
		16#001b# => X"00000000",
		16#001c# => X"00000000",
		16#001d# => X"00000000",
		16#001e# => X"00000000",
		16#001f# => X"00000000",
		16#0020# => X"00000000",
		16#0021# => X"00000000",
		16#0022# => X"00000000",
		16#0023# => X"00000000",
		16#0024# => X"00000000",
		16#0025# => X"00000000",
		16#0026# => X"00000000",
		16#0027# => X"00000000",
		16#0028# => X"00000000",
		16#0029# => X"00000000",
		16#002a# => X"00000000",
		16#002b# => X"00000000",
		16#002c# => X"00000000",
		16#002d# => X"00000000",
		16#002e# => X"00000000",
		16#002f# => X"00000000",
		16#0030# => X"00000000",
		16#0031# => X"00000000",
		16#0032# => X"00000000",
		16#0033# => X"00000000",
		16#0034# => X"00000000",
		16#0035# => X"00000000",
		16#0036# => X"00000000",
		16#0037# => X"00000000",
		16#0038# => X"00000000",
		16#0039# => X"00000000",
		16#003a# => X"00000000",
		16#003b# => X"00000000",
		16#003c# => X"00000000",
		16#003d# => X"00000000",
		16#003e# => X"00000000",
		16#003f# => X"00000000",
		16#0040# => X"18000000",
		16#0041# => X"18200000",
		16#0042# => X"18400000",
		16#0043# => X"18600000",
		16#0044# => X"18800000",
		16#0045# => X"18a00000",
		16#0046# => X"18c00000",
		16#0047# => X"18e00000",
		16#0048# => X"19000000",
		16#0049# => X"19200000",
		16#004a# => X"19400000",
		16#004b# => X"19600000",
		16#004c# => X"19800000",
		16#004d# => X"19a00000",
		16#004e# => X"19c00000",
		16#004f# => X"19e00000",
		16#0050# => X"1a000000",
		16#0051# => X"1a200000",
		16#0052# => X"1a400000",
		16#0053# => X"1a600000",
		16#0054# => X"1a800000",
		16#0055# => X"1aa00000",
		16#0056# => X"1ac00000",
		16#0057# => X"1ae00000",
		16#0058# => X"1b000000",
		16#0059# => X"1b200000",
		16#005a# => X"1b400000",
		16#005b# => X"1b600000",
		16#005c# => X"1b800000",
		16#005d# => X"1ba00000",
		16#005e# => X"1bc00000",
		16#005f# => X"1be00000",
		16#0060# => X"a8200001",
		16#0061# => X"c0000811",
		16#0062# => X"c1400000",
		16#0063# => X"18800000",
		16#0064# => X"a8842028",
		16#0065# => X"44002000",
		16#0066# => X"15000000",
		16#0067# => X"00000000",
		16#0068# => X"00000000",
		16#0069# => X"00000000",
		16#006a# => X"00000000",
		16#006b# => X"00000000",
		16#006c# => X"00000000",
		16#006d# => X"00000000",
		16#006e# => X"00000000",
		16#006f# => X"00000000",
		16#0070# => X"00000000",
		16#0071# => X"00000000",
		16#0072# => X"00000000",
		16#0073# => X"00000000",
		16#0074# => X"00000000",
		16#0075# => X"00000000",
		16#0076# => X"00000000",
		16#0077# => X"00000000",
		16#0078# => X"00000000",
		16#0079# => X"00000000",
		16#007a# => X"00000000",
		16#007b# => X"00000000",
		16#007c# => X"00000000",
		16#007d# => X"00000000",
		16#007e# => X"00000000",
		16#007f# => X"00000000",
		16#0080# => X"9c21ff00",
		16#0081# => X"d4011804",
		16#0082# => X"d4012008",
		16#0083# => X"b4600010",
		16#0084# => X"00003424",
		16#0085# => X"b4800020",
		16#0086# => X"00000000",
		16#0087# => X"00000000",
		16#0088# => X"00000000",
		16#0089# => X"00000000",
		16#008a# => X"00000000",
		16#008b# => X"00000000",
		16#008c# => X"00000000",
		16#008d# => X"00000000",
		16#008e# => X"00000000",
		16#008f# => X"00000000",
		16#0090# => X"00000000",
		16#0091# => X"00000000",
		16#0092# => X"00000000",
		16#0093# => X"00000000",
		16#0094# => X"00000000",
		16#0095# => X"00000000",
		16#0096# => X"00000000",
		16#0097# => X"00000000",
		16#0098# => X"00000000",
		16#0099# => X"00000000",
		16#009a# => X"00000000",
		16#009b# => X"00000000",
		16#009c# => X"00000000",
		16#009d# => X"00000000",
		16#009e# => X"00000000",
		16#009f# => X"00000000",
		16#00a0# => X"00000000",
		16#00a1# => X"00000000",
		16#00a2# => X"00000000",
		16#00a3# => X"00000000",
		16#00a4# => X"00000000",
		16#00a5# => X"00000000",
		16#00a6# => X"00000000",
		16#00a7# => X"00000000",
		16#00a8# => X"00000000",
		16#00a9# => X"00000000",
		16#00aa# => X"00000000",
		16#00ab# => X"00000000",
		16#00ac# => X"00000000",
		16#00ad# => X"00000000",
		16#00ae# => X"00000000",
		16#00af# => X"00000000",
		16#00b0# => X"00000000",
		16#00b1# => X"00000000",
		16#00b2# => X"00000000",
		16#00b3# => X"00000000",
		16#00b4# => X"00000000",
		16#00b5# => X"00000000",
		16#00b6# => X"00000000",
		16#00b7# => X"00000000",
		16#00b8# => X"00000000",
		16#00b9# => X"00000000",
		16#00ba# => X"00000000",
		16#00bb# => X"00000000",
		16#00bc# => X"00000000",
		16#00bd# => X"00000000",
		16#00be# => X"00000000",
		16#00bf# => X"00000000",
		16#00c0# => X"9c21ff00",
		16#00c1# => X"d4011804",
		16#00c2# => X"d4012008",
		16#00c3# => X"b4600010",
		16#00c4# => X"000033e4",
		16#00c5# => X"b4800020",
		16#00c6# => X"00000000",
		16#00c7# => X"00000000",
		16#00c8# => X"00000000",
		16#00c9# => X"00000000",
		16#00ca# => X"00000000",
		16#00cb# => X"00000000",
		16#00cc# => X"00000000",
		16#00cd# => X"00000000",
		16#00ce# => X"00000000",
		16#00cf# => X"00000000",
		16#00d0# => X"00000000",
		16#00d1# => X"00000000",
		16#00d2# => X"00000000",
		16#00d3# => X"00000000",
		16#00d4# => X"00000000",
		16#00d5# => X"00000000",
		16#00d6# => X"00000000",
		16#00d7# => X"00000000",
		16#00d8# => X"00000000",
		16#00d9# => X"00000000",
		16#00da# => X"00000000",
		16#00db# => X"00000000",
		16#00dc# => X"00000000",
		16#00dd# => X"00000000",
		16#00de# => X"00000000",
		16#00df# => X"00000000",
		16#00e0# => X"00000000",
		16#00e1# => X"00000000",
		16#00e2# => X"00000000",
		16#00e3# => X"00000000",
		16#00e4# => X"00000000",
		16#00e5# => X"00000000",
		16#00e6# => X"00000000",
		16#00e7# => X"00000000",
		16#00e8# => X"00000000",
		16#00e9# => X"00000000",
		16#00ea# => X"00000000",
		16#00eb# => X"00000000",
		16#00ec# => X"00000000",
		16#00ed# => X"00000000",
		16#00ee# => X"00000000",
		16#00ef# => X"00000000",
		16#00f0# => X"00000000",
		16#00f1# => X"00000000",
		16#00f2# => X"00000000",
		16#00f3# => X"00000000",
		16#00f4# => X"00000000",
		16#00f5# => X"00000000",
		16#00f6# => X"00000000",
		16#00f7# => X"00000000",
		16#00f8# => X"00000000",
		16#00f9# => X"00000000",
		16#00fa# => X"00000000",
		16#00fb# => X"00000000",
		16#00fc# => X"00000000",
		16#00fd# => X"00000000",
		16#00fe# => X"00000000",
		16#00ff# => X"00000000",
		16#0100# => X"9c21ff00",
		16#0101# => X"d4011804",
		16#0102# => X"d4012008",
		16#0103# => X"b4600010",
		16#0104# => X"000033a4",
		16#0105# => X"b4800020",
		16#0106# => X"00000000",
		16#0107# => X"00000000",
		16#0108# => X"00000000",
		16#0109# => X"00000000",
		16#010a# => X"00000000",
		16#010b# => X"00000000",
		16#010c# => X"00000000",
		16#010d# => X"00000000",
		16#010e# => X"00000000",
		16#010f# => X"00000000",
		16#0110# => X"00000000",
		16#0111# => X"00000000",
		16#0112# => X"00000000",
		16#0113# => X"00000000",
		16#0114# => X"00000000",
		16#0115# => X"00000000",
		16#0116# => X"00000000",
		16#0117# => X"00000000",
		16#0118# => X"00000000",
		16#0119# => X"00000000",
		16#011a# => X"00000000",
		16#011b# => X"00000000",
		16#011c# => X"00000000",
		16#011d# => X"00000000",
		16#011e# => X"00000000",
		16#011f# => X"00000000",
		16#0120# => X"00000000",
		16#0121# => X"00000000",
		16#0122# => X"00000000",
		16#0123# => X"00000000",
		16#0124# => X"00000000",
		16#0125# => X"00000000",
		16#0126# => X"00000000",
		16#0127# => X"00000000",
		16#0128# => X"00000000",
		16#0129# => X"00000000",
		16#012a# => X"00000000",
		16#012b# => X"00000000",
		16#012c# => X"00000000",
		16#012d# => X"00000000",
		16#012e# => X"00000000",
		16#012f# => X"00000000",
		16#0130# => X"00000000",
		16#0131# => X"00000000",
		16#0132# => X"00000000",
		16#0133# => X"00000000",
		16#0134# => X"00000000",
		16#0135# => X"00000000",
		16#0136# => X"00000000",
		16#0137# => X"00000000",
		16#0138# => X"00000000",
		16#0139# => X"00000000",
		16#013a# => X"00000000",
		16#013b# => X"00000000",
		16#013c# => X"00000000",
		16#013d# => X"00000000",
		16#013e# => X"00000000",
		16#013f# => X"00000000",
		16#0140# => X"9c21ff00",
		16#0141# => X"d4011804",
		16#0142# => X"d4012008",
		16#0143# => X"b4600010",
		16#0144# => X"00003364",
		16#0145# => X"b4800020",
		16#0146# => X"00000000",
		16#0147# => X"00000000",
		16#0148# => X"00000000",
		16#0149# => X"00000000",
		16#014a# => X"00000000",
		16#014b# => X"00000000",
		16#014c# => X"00000000",
		16#014d# => X"00000000",
		16#014e# => X"00000000",
		16#014f# => X"00000000",
		16#0150# => X"00000000",
		16#0151# => X"00000000",
		16#0152# => X"00000000",
		16#0153# => X"00000000",
		16#0154# => X"00000000",
		16#0155# => X"00000000",
		16#0156# => X"00000000",
		16#0157# => X"00000000",
		16#0158# => X"00000000",
		16#0159# => X"00000000",
		16#015a# => X"00000000",
		16#015b# => X"00000000",
		16#015c# => X"00000000",
		16#015d# => X"00000000",
		16#015e# => X"00000000",
		16#015f# => X"00000000",
		16#0160# => X"00000000",
		16#0161# => X"00000000",
		16#0162# => X"00000000",
		16#0163# => X"00000000",
		16#0164# => X"00000000",
		16#0165# => X"00000000",
		16#0166# => X"00000000",
		16#0167# => X"00000000",
		16#0168# => X"00000000",
		16#0169# => X"00000000",
		16#016a# => X"00000000",
		16#016b# => X"00000000",
		16#016c# => X"00000000",
		16#016d# => X"00000000",
		16#016e# => X"00000000",
		16#016f# => X"00000000",
		16#0170# => X"00000000",
		16#0171# => X"00000000",
		16#0172# => X"00000000",
		16#0173# => X"00000000",
		16#0174# => X"00000000",
		16#0175# => X"00000000",
		16#0176# => X"00000000",
		16#0177# => X"00000000",
		16#0178# => X"00000000",
		16#0179# => X"00000000",
		16#017a# => X"00000000",
		16#017b# => X"00000000",
		16#017c# => X"00000000",
		16#017d# => X"00000000",
		16#017e# => X"00000000",
		16#017f# => X"00000000",
		16#0180# => X"9c21ff00",
		16#0181# => X"d4011804",
		16#0182# => X"d4012008",
		16#0183# => X"b4600010",
		16#0184# => X"00003324",
		16#0185# => X"b4800020",
		16#0186# => X"00000000",
		16#0187# => X"00000000",
		16#0188# => X"00000000",
		16#0189# => X"00000000",
		16#018a# => X"00000000",
		16#018b# => X"00000000",
		16#018c# => X"00000000",
		16#018d# => X"00000000",
		16#018e# => X"00000000",
		16#018f# => X"00000000",
		16#0190# => X"00000000",
		16#0191# => X"00000000",
		16#0192# => X"00000000",
		16#0193# => X"00000000",
		16#0194# => X"00000000",
		16#0195# => X"00000000",
		16#0196# => X"00000000",
		16#0197# => X"00000000",
		16#0198# => X"00000000",
		16#0199# => X"00000000",
		16#019a# => X"00000000",
		16#019b# => X"00000000",
		16#019c# => X"00000000",
		16#019d# => X"00000000",
		16#019e# => X"00000000",
		16#019f# => X"00000000",
		16#01a0# => X"00000000",
		16#01a1# => X"00000000",
		16#01a2# => X"00000000",
		16#01a3# => X"00000000",
		16#01a4# => X"00000000",
		16#01a5# => X"00000000",
		16#01a6# => X"00000000",
		16#01a7# => X"00000000",
		16#01a8# => X"00000000",
		16#01a9# => X"00000000",
		16#01aa# => X"00000000",
		16#01ab# => X"00000000",
		16#01ac# => X"00000000",
		16#01ad# => X"00000000",
		16#01ae# => X"00000000",
		16#01af# => X"00000000",
		16#01b0# => X"00000000",
		16#01b1# => X"00000000",
		16#01b2# => X"00000000",
		16#01b3# => X"00000000",
		16#01b4# => X"00000000",
		16#01b5# => X"00000000",
		16#01b6# => X"00000000",
		16#01b7# => X"00000000",
		16#01b8# => X"00000000",
		16#01b9# => X"00000000",
		16#01ba# => X"00000000",
		16#01bb# => X"00000000",
		16#01bc# => X"00000000",
		16#01bd# => X"00000000",
		16#01be# => X"00000000",
		16#01bf# => X"00000000",
		16#01c0# => X"9c21ff00",
		16#01c1# => X"d4011804",
		16#01c2# => X"d4012008",
		16#01c3# => X"b4600010",
		16#01c4# => X"000032e4",
		16#01c5# => X"b4800020",
		16#01c6# => X"00000000",
		16#01c7# => X"00000000",
		16#01c8# => X"00000000",
		16#01c9# => X"00000000",
		16#01ca# => X"00000000",
		16#01cb# => X"00000000",
		16#01cc# => X"00000000",
		16#01cd# => X"00000000",
		16#01ce# => X"00000000",
		16#01cf# => X"00000000",
		16#01d0# => X"00000000",
		16#01d1# => X"00000000",
		16#01d2# => X"00000000",
		16#01d3# => X"00000000",
		16#01d4# => X"00000000",
		16#01d5# => X"00000000",
		16#01d6# => X"00000000",
		16#01d7# => X"00000000",
		16#01d8# => X"00000000",
		16#01d9# => X"00000000",
		16#01da# => X"00000000",
		16#01db# => X"00000000",
		16#01dc# => X"00000000",
		16#01dd# => X"00000000",
		16#01de# => X"00000000",
		16#01df# => X"00000000",
		16#01e0# => X"00000000",
		16#01e1# => X"00000000",
		16#01e2# => X"00000000",
		16#01e3# => X"00000000",
		16#01e4# => X"00000000",
		16#01e5# => X"00000000",
		16#01e6# => X"00000000",
		16#01e7# => X"00000000",
		16#01e8# => X"00000000",
		16#01e9# => X"00000000",
		16#01ea# => X"00000000",
		16#01eb# => X"00000000",
		16#01ec# => X"00000000",
		16#01ed# => X"00000000",
		16#01ee# => X"00000000",
		16#01ef# => X"00000000",
		16#01f0# => X"00000000",
		16#01f1# => X"00000000",
		16#01f2# => X"00000000",
		16#01f3# => X"00000000",
		16#01f4# => X"00000000",
		16#01f5# => X"00000000",
		16#01f6# => X"00000000",
		16#01f7# => X"00000000",
		16#01f8# => X"00000000",
		16#01f9# => X"00000000",
		16#01fa# => X"00000000",
		16#01fb# => X"00000000",
		16#01fc# => X"00000000",
		16#01fd# => X"00000000",
		16#01fe# => X"00000000",
		16#01ff# => X"00000000",
		16#0200# => X"9c21ff00",
		16#0201# => X"d4011804",
		16#0202# => X"d4012008",
		16#0203# => X"b4600010",
		16#0204# => X"000032a4",
		16#0205# => X"b4800020",
		16#0206# => X"00000000",
		16#0207# => X"00000000",
		16#0208# => X"00000000",
		16#0209# => X"00000000",
		16#020a# => X"00000000",
		16#020b# => X"00000000",
		16#020c# => X"00000000",
		16#020d# => X"00000000",
		16#020e# => X"00000000",
		16#020f# => X"00000000",
		16#0210# => X"00000000",
		16#0211# => X"00000000",
		16#0212# => X"00000000",
		16#0213# => X"00000000",
		16#0214# => X"00000000",
		16#0215# => X"00000000",
		16#0216# => X"00000000",
		16#0217# => X"00000000",
		16#0218# => X"00000000",
		16#0219# => X"00000000",
		16#021a# => X"00000000",
		16#021b# => X"00000000",
		16#021c# => X"00000000",
		16#021d# => X"00000000",
		16#021e# => X"00000000",
		16#021f# => X"00000000",
		16#0220# => X"00000000",
		16#0221# => X"00000000",
		16#0222# => X"00000000",
		16#0223# => X"00000000",
		16#0224# => X"00000000",
		16#0225# => X"00000000",
		16#0226# => X"00000000",
		16#0227# => X"00000000",
		16#0228# => X"00000000",
		16#0229# => X"00000000",
		16#022a# => X"00000000",
		16#022b# => X"00000000",
		16#022c# => X"00000000",
		16#022d# => X"00000000",
		16#022e# => X"00000000",
		16#022f# => X"00000000",
		16#0230# => X"00000000",
		16#0231# => X"00000000",
		16#0232# => X"00000000",
		16#0233# => X"00000000",
		16#0234# => X"00000000",
		16#0235# => X"00000000",
		16#0236# => X"00000000",
		16#0237# => X"00000000",
		16#0238# => X"00000000",
		16#0239# => X"00000000",
		16#023a# => X"00000000",
		16#023b# => X"00000000",
		16#023c# => X"00000000",
		16#023d# => X"00000000",
		16#023e# => X"00000000",
		16#023f# => X"00000000",
		16#0240# => X"9c21ff00",
		16#0241# => X"d4011804",
		16#0242# => X"d4012008",
		16#0243# => X"b4600010",
		16#0244# => X"00003264",
		16#0245# => X"b4800020",
		16#0246# => X"00000000",
		16#0247# => X"00000000",
		16#0248# => X"00000000",
		16#0249# => X"00000000",
		16#024a# => X"00000000",
		16#024b# => X"00000000",
		16#024c# => X"00000000",
		16#024d# => X"00000000",
		16#024e# => X"00000000",
		16#024f# => X"00000000",
		16#0250# => X"00000000",
		16#0251# => X"00000000",
		16#0252# => X"00000000",
		16#0253# => X"00000000",
		16#0254# => X"00000000",
		16#0255# => X"00000000",
		16#0256# => X"00000000",
		16#0257# => X"00000000",
		16#0258# => X"00000000",
		16#0259# => X"00000000",
		16#025a# => X"00000000",
		16#025b# => X"00000000",
		16#025c# => X"00000000",
		16#025d# => X"00000000",
		16#025e# => X"00000000",
		16#025f# => X"00000000",
		16#0260# => X"00000000",
		16#0261# => X"00000000",
		16#0262# => X"00000000",
		16#0263# => X"00000000",
		16#0264# => X"00000000",
		16#0265# => X"00000000",
		16#0266# => X"00000000",
		16#0267# => X"00000000",
		16#0268# => X"00000000",
		16#0269# => X"00000000",
		16#026a# => X"00000000",
		16#026b# => X"00000000",
		16#026c# => X"00000000",
		16#026d# => X"00000000",
		16#026e# => X"00000000",
		16#026f# => X"00000000",
		16#0270# => X"00000000",
		16#0271# => X"00000000",
		16#0272# => X"00000000",
		16#0273# => X"00000000",
		16#0274# => X"00000000",
		16#0275# => X"00000000",
		16#0276# => X"00000000",
		16#0277# => X"00000000",
		16#0278# => X"00000000",
		16#0279# => X"00000000",
		16#027a# => X"00000000",
		16#027b# => X"00000000",
		16#027c# => X"00000000",
		16#027d# => X"00000000",
		16#027e# => X"00000000",
		16#027f# => X"00000000",
		16#0280# => X"9c21ff00",
		16#0281# => X"d4011804",
		16#0282# => X"d4012008",
		16#0283# => X"b4600010",
		16#0284# => X"00003224",
		16#0285# => X"b4800020",
		16#0286# => X"00000000",
		16#0287# => X"00000000",
		16#0288# => X"00000000",
		16#0289# => X"00000000",
		16#028a# => X"00000000",
		16#028b# => X"00000000",
		16#028c# => X"00000000",
		16#028d# => X"00000000",
		16#028e# => X"00000000",
		16#028f# => X"00000000",
		16#0290# => X"00000000",
		16#0291# => X"00000000",
		16#0292# => X"00000000",
		16#0293# => X"00000000",
		16#0294# => X"00000000",
		16#0295# => X"00000000",
		16#0296# => X"00000000",
		16#0297# => X"00000000",
		16#0298# => X"00000000",
		16#0299# => X"00000000",
		16#029a# => X"00000000",
		16#029b# => X"00000000",
		16#029c# => X"00000000",
		16#029d# => X"00000000",
		16#029e# => X"00000000",
		16#029f# => X"00000000",
		16#02a0# => X"00000000",
		16#02a1# => X"00000000",
		16#02a2# => X"00000000",
		16#02a3# => X"00000000",
		16#02a4# => X"00000000",
		16#02a5# => X"00000000",
		16#02a6# => X"00000000",
		16#02a7# => X"00000000",
		16#02a8# => X"00000000",
		16#02a9# => X"00000000",
		16#02aa# => X"00000000",
		16#02ab# => X"00000000",
		16#02ac# => X"00000000",
		16#02ad# => X"00000000",
		16#02ae# => X"00000000",
		16#02af# => X"00000000",
		16#02b0# => X"00000000",
		16#02b1# => X"00000000",
		16#02b2# => X"00000000",
		16#02b3# => X"00000000",
		16#02b4# => X"00000000",
		16#02b5# => X"00000000",
		16#02b6# => X"00000000",
		16#02b7# => X"00000000",
		16#02b8# => X"00000000",
		16#02b9# => X"00000000",
		16#02ba# => X"00000000",
		16#02bb# => X"00000000",
		16#02bc# => X"00000000",
		16#02bd# => X"00000000",
		16#02be# => X"00000000",
		16#02bf# => X"00000000",
		16#02c0# => X"9c21ff00",
		16#02c1# => X"d4011804",
		16#02c2# => X"d4012008",
		16#02c3# => X"b4600010",
		16#02c4# => X"000031e4",
		16#02c5# => X"b4800020",
		16#02c6# => X"00000000",
		16#02c7# => X"00000000",
		16#02c8# => X"00000000",
		16#02c9# => X"00000000",
		16#02ca# => X"00000000",
		16#02cb# => X"00000000",
		16#02cc# => X"00000000",
		16#02cd# => X"00000000",
		16#02ce# => X"00000000",
		16#02cf# => X"00000000",
		16#02d0# => X"00000000",
		16#02d1# => X"00000000",
		16#02d2# => X"00000000",
		16#02d3# => X"00000000",
		16#02d4# => X"00000000",
		16#02d5# => X"00000000",
		16#02d6# => X"00000000",
		16#02d7# => X"00000000",
		16#02d8# => X"00000000",
		16#02d9# => X"00000000",
		16#02da# => X"00000000",
		16#02db# => X"00000000",
		16#02dc# => X"00000000",
		16#02dd# => X"00000000",
		16#02de# => X"00000000",
		16#02df# => X"00000000",
		16#02e0# => X"00000000",
		16#02e1# => X"00000000",
		16#02e2# => X"00000000",
		16#02e3# => X"00000000",
		16#02e4# => X"00000000",
		16#02e5# => X"00000000",
		16#02e6# => X"00000000",
		16#02e7# => X"00000000",
		16#02e8# => X"00000000",
		16#02e9# => X"00000000",
		16#02ea# => X"00000000",
		16#02eb# => X"00000000",
		16#02ec# => X"00000000",
		16#02ed# => X"00000000",
		16#02ee# => X"00000000",
		16#02ef# => X"00000000",
		16#02f0# => X"00000000",
		16#02f1# => X"00000000",
		16#02f2# => X"00000000",
		16#02f3# => X"00000000",
		16#02f4# => X"00000000",
		16#02f5# => X"00000000",
		16#02f6# => X"00000000",
		16#02f7# => X"00000000",
		16#02f8# => X"00000000",
		16#02f9# => X"00000000",
		16#02fa# => X"00000000",
		16#02fb# => X"00000000",
		16#02fc# => X"00000000",
		16#02fd# => X"00000000",
		16#02fe# => X"00000000",
		16#02ff# => X"00000000",
		16#0300# => X"9c21ff00",
		16#0301# => X"d4011804",
		16#0302# => X"d4012008",
		16#0303# => X"b4600010",
		16#0304# => X"000031a4",
		16#0305# => X"b4800020",
		16#0306# => X"00000000",
		16#0307# => X"00000000",
		16#0308# => X"00000000",
		16#0309# => X"00000000",
		16#030a# => X"00000000",
		16#030b# => X"00000000",
		16#030c# => X"00000000",
		16#030d# => X"00000000",
		16#030e# => X"00000000",
		16#030f# => X"00000000",
		16#0310# => X"00000000",
		16#0311# => X"00000000",
		16#0312# => X"00000000",
		16#0313# => X"00000000",
		16#0314# => X"00000000",
		16#0315# => X"00000000",
		16#0316# => X"00000000",
		16#0317# => X"00000000",
		16#0318# => X"00000000",
		16#0319# => X"00000000",
		16#031a# => X"00000000",
		16#031b# => X"00000000",
		16#031c# => X"00000000",
		16#031d# => X"00000000",
		16#031e# => X"00000000",
		16#031f# => X"00000000",
		16#0320# => X"00000000",
		16#0321# => X"00000000",
		16#0322# => X"00000000",
		16#0323# => X"00000000",
		16#0324# => X"00000000",
		16#0325# => X"00000000",
		16#0326# => X"00000000",
		16#0327# => X"00000000",
		16#0328# => X"00000000",
		16#0329# => X"00000000",
		16#032a# => X"00000000",
		16#032b# => X"00000000",
		16#032c# => X"00000000",
		16#032d# => X"00000000",
		16#032e# => X"00000000",
		16#032f# => X"00000000",
		16#0330# => X"00000000",
		16#0331# => X"00000000",
		16#0332# => X"00000000",
		16#0333# => X"00000000",
		16#0334# => X"00000000",
		16#0335# => X"00000000",
		16#0336# => X"00000000",
		16#0337# => X"00000000",
		16#0338# => X"00000000",
		16#0339# => X"00000000",
		16#033a# => X"00000000",
		16#033b# => X"00000000",
		16#033c# => X"00000000",
		16#033d# => X"00000000",
		16#033e# => X"00000000",
		16#033f# => X"00000000",
		16#0340# => X"9c21ff00",
		16#0341# => X"d4011804",
		16#0342# => X"d4012008",
		16#0343# => X"b4600010",
		16#0344# => X"00003164",
		16#0345# => X"b4800020",
		16#0346# => X"00000000",
		16#0347# => X"00000000",
		16#0348# => X"00000000",
		16#0349# => X"00000000",
		16#034a# => X"00000000",
		16#034b# => X"00000000",
		16#034c# => X"00000000",
		16#034d# => X"00000000",
		16#034e# => X"00000000",
		16#034f# => X"00000000",
		16#0350# => X"00000000",
		16#0351# => X"00000000",
		16#0352# => X"00000000",
		16#0353# => X"00000000",
		16#0354# => X"00000000",
		16#0355# => X"00000000",
		16#0356# => X"00000000",
		16#0357# => X"00000000",
		16#0358# => X"00000000",
		16#0359# => X"00000000",
		16#035a# => X"00000000",
		16#035b# => X"00000000",
		16#035c# => X"00000000",
		16#035d# => X"00000000",
		16#035e# => X"00000000",
		16#035f# => X"00000000",
		16#0360# => X"00000000",
		16#0361# => X"00000000",
		16#0362# => X"00000000",
		16#0363# => X"00000000",
		16#0364# => X"00000000",
		16#0365# => X"00000000",
		16#0366# => X"00000000",
		16#0367# => X"00000000",
		16#0368# => X"00000000",
		16#0369# => X"00000000",
		16#036a# => X"00000000",
		16#036b# => X"00000000",
		16#036c# => X"00000000",
		16#036d# => X"00000000",
		16#036e# => X"00000000",
		16#036f# => X"00000000",
		16#0370# => X"00000000",
		16#0371# => X"00000000",
		16#0372# => X"00000000",
		16#0373# => X"00000000",
		16#0374# => X"00000000",
		16#0375# => X"00000000",
		16#0376# => X"00000000",
		16#0377# => X"00000000",
		16#0378# => X"00000000",
		16#0379# => X"00000000",
		16#037a# => X"00000000",
		16#037b# => X"00000000",
		16#037c# => X"00000000",
		16#037d# => X"00000000",
		16#037e# => X"00000000",
		16#037f# => X"00000000",
		16#0380# => X"9c21ff00",
		16#0381# => X"d4011804",
		16#0382# => X"d4012008",
		16#0383# => X"b4600010",
		16#0384# => X"00003124",
		16#0385# => X"b4800020",
		16#0386# => X"00000000",
		16#0387# => X"00000000",
		16#0388# => X"00000000",
		16#0389# => X"00000000",
		16#038a# => X"00000000",
		16#038b# => X"00000000",
		16#038c# => X"00000000",
		16#038d# => X"00000000",
		16#038e# => X"00000000",
		16#038f# => X"00000000",
		16#0390# => X"00000000",
		16#0391# => X"00000000",
		16#0392# => X"00000000",
		16#0393# => X"00000000",
		16#0394# => X"00000000",
		16#0395# => X"00000000",
		16#0396# => X"00000000",
		16#0397# => X"00000000",
		16#0398# => X"00000000",
		16#0399# => X"00000000",
		16#039a# => X"00000000",
		16#039b# => X"00000000",
		16#039c# => X"00000000",
		16#039d# => X"00000000",
		16#039e# => X"00000000",
		16#039f# => X"00000000",
		16#03a0# => X"00000000",
		16#03a1# => X"00000000",
		16#03a2# => X"00000000",
		16#03a3# => X"00000000",
		16#03a4# => X"00000000",
		16#03a5# => X"00000000",
		16#03a6# => X"00000000",
		16#03a7# => X"00000000",
		16#03a8# => X"00000000",
		16#03a9# => X"00000000",
		16#03aa# => X"00000000",
		16#03ab# => X"00000000",
		16#03ac# => X"00000000",
		16#03ad# => X"00000000",
		16#03ae# => X"00000000",
		16#03af# => X"00000000",
		16#03b0# => X"00000000",
		16#03b1# => X"00000000",
		16#03b2# => X"00000000",
		16#03b3# => X"00000000",
		16#03b4# => X"00000000",
		16#03b5# => X"00000000",
		16#03b6# => X"00000000",
		16#03b7# => X"00000000",
		16#03b8# => X"00000000",
		16#03b9# => X"00000000",
		16#03ba# => X"00000000",
		16#03bb# => X"00000000",
		16#03bc# => X"00000000",
		16#03bd# => X"00000000",
		16#03be# => X"00000000",
		16#03bf# => X"00000000",
		16#03c0# => X"9c21ff00",
		16#03c1# => X"d4011804",
		16#03c2# => X"d4012008",
		16#03c3# => X"b4600010",
		16#03c4# => X"000030e4",
		16#03c5# => X"b4800020",
		16#03c6# => X"00000000",
		16#03c7# => X"00000000",
		16#03c8# => X"00000000",
		16#03c9# => X"00000000",
		16#03ca# => X"00000000",
		16#03cb# => X"00000000",
		16#03cc# => X"00000000",
		16#03cd# => X"00000000",
		16#03ce# => X"00000000",
		16#03cf# => X"00000000",
		16#03d0# => X"00000000",
		16#03d1# => X"00000000",
		16#03d2# => X"00000000",
		16#03d3# => X"00000000",
		16#03d4# => X"00000000",
		16#03d5# => X"00000000",
		16#03d6# => X"00000000",
		16#03d7# => X"00000000",
		16#03d8# => X"00000000",
		16#03d9# => X"00000000",
		16#03da# => X"00000000",
		16#03db# => X"00000000",
		16#03dc# => X"00000000",
		16#03dd# => X"00000000",
		16#03de# => X"00000000",
		16#03df# => X"00000000",
		16#03e0# => X"00000000",
		16#03e1# => X"00000000",
		16#03e2# => X"00000000",
		16#03e3# => X"00000000",
		16#03e4# => X"00000000",
		16#03e5# => X"00000000",
		16#03e6# => X"00000000",
		16#03e7# => X"00000000",
		16#03e8# => X"00000000",
		16#03e9# => X"00000000",
		16#03ea# => X"00000000",
		16#03eb# => X"00000000",
		16#03ec# => X"00000000",
		16#03ed# => X"00000000",
		16#03ee# => X"00000000",
		16#03ef# => X"00000000",
		16#03f0# => X"00000000",
		16#03f1# => X"00000000",
		16#03f2# => X"00000000",
		16#03f3# => X"00000000",
		16#03f4# => X"00000000",
		16#03f5# => X"00000000",
		16#03f6# => X"00000000",
		16#03f7# => X"00000000",
		16#03f8# => X"00000000",
		16#03f9# => X"00000000",
		16#03fa# => X"00000000",
		16#03fb# => X"00000000",
		16#03fc# => X"00000000",
		16#03fd# => X"00000000",
		16#03fe# => X"00000000",
		16#03ff# => X"00000000",
		16#0400# => X"9c21ff00",
		16#0401# => X"d4011804",
		16#0402# => X"d4012008",
		16#0403# => X"b4600010",
		16#0404# => X"000030a4",
		16#0405# => X"b4800020",
		16#0406# => X"00000000",
		16#0407# => X"00000000",
		16#0408# => X"00000000",
		16#0409# => X"00000000",
		16#040a# => X"00000000",
		16#040b# => X"00000000",
		16#040c# => X"00000000",
		16#040d# => X"00000000",
		16#040e# => X"00000000",
		16#040f# => X"00000000",
		16#0410# => X"00000000",
		16#0411# => X"00000000",
		16#0412# => X"00000000",
		16#0413# => X"00000000",
		16#0414# => X"00000000",
		16#0415# => X"00000000",
		16#0416# => X"00000000",
		16#0417# => X"00000000",
		16#0418# => X"00000000",
		16#0419# => X"00000000",
		16#041a# => X"00000000",
		16#041b# => X"00000000",
		16#041c# => X"00000000",
		16#041d# => X"00000000",
		16#041e# => X"00000000",
		16#041f# => X"00000000",
		16#0420# => X"00000000",
		16#0421# => X"00000000",
		16#0422# => X"00000000",
		16#0423# => X"00000000",
		16#0424# => X"00000000",
		16#0425# => X"00000000",
		16#0426# => X"00000000",
		16#0427# => X"00000000",
		16#0428# => X"00000000",
		16#0429# => X"00000000",
		16#042a# => X"00000000",
		16#042b# => X"00000000",
		16#042c# => X"00000000",
		16#042d# => X"00000000",
		16#042e# => X"00000000",
		16#042f# => X"00000000",
		16#0430# => X"00000000",
		16#0431# => X"00000000",
		16#0432# => X"00000000",
		16#0433# => X"00000000",
		16#0434# => X"00000000",
		16#0435# => X"00000000",
		16#0436# => X"00000000",
		16#0437# => X"00000000",
		16#0438# => X"00000000",
		16#0439# => X"00000000",
		16#043a# => X"00000000",
		16#043b# => X"00000000",
		16#043c# => X"00000000",
		16#043d# => X"00000000",
		16#043e# => X"00000000",
		16#043f# => X"00000000",
		16#0440# => X"9c21ff00",
		16#0441# => X"d4011804",
		16#0442# => X"d4012008",
		16#0443# => X"b4600010",
		16#0444# => X"00003064",
		16#0445# => X"b4800020",
		16#0446# => X"00000000",
		16#0447# => X"00000000",
		16#0448# => X"00000000",
		16#0449# => X"00000000",
		16#044a# => X"00000000",
		16#044b# => X"00000000",
		16#044c# => X"00000000",
		16#044d# => X"00000000",
		16#044e# => X"00000000",
		16#044f# => X"00000000",
		16#0450# => X"00000000",
		16#0451# => X"00000000",
		16#0452# => X"00000000",
		16#0453# => X"00000000",
		16#0454# => X"00000000",
		16#0455# => X"00000000",
		16#0456# => X"00000000",
		16#0457# => X"00000000",
		16#0458# => X"00000000",
		16#0459# => X"00000000",
		16#045a# => X"00000000",
		16#045b# => X"00000000",
		16#045c# => X"00000000",
		16#045d# => X"00000000",
		16#045e# => X"00000000",
		16#045f# => X"00000000",
		16#0460# => X"00000000",
		16#0461# => X"00000000",
		16#0462# => X"00000000",
		16#0463# => X"00000000",
		16#0464# => X"00000000",
		16#0465# => X"00000000",
		16#0466# => X"00000000",
		16#0467# => X"00000000",
		16#0468# => X"00000000",
		16#0469# => X"00000000",
		16#046a# => X"00000000",
		16#046b# => X"00000000",
		16#046c# => X"00000000",
		16#046d# => X"00000000",
		16#046e# => X"00000000",
		16#046f# => X"00000000",
		16#0470# => X"00000000",
		16#0471# => X"00000000",
		16#0472# => X"00000000",
		16#0473# => X"00000000",
		16#0474# => X"00000000",
		16#0475# => X"00000000",
		16#0476# => X"00000000",
		16#0477# => X"00000000",
		16#0478# => X"00000000",
		16#0479# => X"00000000",
		16#047a# => X"00000000",
		16#047b# => X"00000000",
		16#047c# => X"00000000",
		16#047d# => X"00000000",
		16#047e# => X"00000000",
		16#047f# => X"00000000",
		16#0480# => X"9c21ff00",
		16#0481# => X"d4011804",
		16#0482# => X"d4012008",
		16#0483# => X"b4600010",
		16#0484# => X"00003024",
		16#0485# => X"b4800020",
		16#0486# => X"00000000",
		16#0487# => X"00000000",
		16#0488# => X"00000000",
		16#0489# => X"00000000",
		16#048a# => X"00000000",
		16#048b# => X"00000000",
		16#048c# => X"00000000",
		16#048d# => X"00000000",
		16#048e# => X"00000000",
		16#048f# => X"00000000",
		16#0490# => X"00000000",
		16#0491# => X"00000000",
		16#0492# => X"00000000",
		16#0493# => X"00000000",
		16#0494# => X"00000000",
		16#0495# => X"00000000",
		16#0496# => X"00000000",
		16#0497# => X"00000000",
		16#0498# => X"00000000",
		16#0499# => X"00000000",
		16#049a# => X"00000000",
		16#049b# => X"00000000",
		16#049c# => X"00000000",
		16#049d# => X"00000000",
		16#049e# => X"00000000",
		16#049f# => X"00000000",
		16#04a0# => X"00000000",
		16#04a1# => X"00000000",
		16#04a2# => X"00000000",
		16#04a3# => X"00000000",
		16#04a4# => X"00000000",
		16#04a5# => X"00000000",
		16#04a6# => X"00000000",
		16#04a7# => X"00000000",
		16#04a8# => X"00000000",
		16#04a9# => X"00000000",
		16#04aa# => X"00000000",
		16#04ab# => X"00000000",
		16#04ac# => X"00000000",
		16#04ad# => X"00000000",
		16#04ae# => X"00000000",
		16#04af# => X"00000000",
		16#04b0# => X"00000000",
		16#04b1# => X"00000000",
		16#04b2# => X"00000000",
		16#04b3# => X"00000000",
		16#04b4# => X"00000000",
		16#04b5# => X"00000000",
		16#04b6# => X"00000000",
		16#04b7# => X"00000000",
		16#04b8# => X"00000000",
		16#04b9# => X"00000000",
		16#04ba# => X"00000000",
		16#04bb# => X"00000000",
		16#04bc# => X"00000000",
		16#04bd# => X"00000000",
		16#04be# => X"00000000",
		16#04bf# => X"00000000",
		16#04c0# => X"9c21ff00",
		16#04c1# => X"d4011804",
		16#04c2# => X"d4012008",
		16#04c3# => X"b4600010",
		16#04c4# => X"00002fe4",
		16#04c5# => X"b4800020",
		16#04c6# => X"00000000",
		16#04c7# => X"00000000",
		16#04c8# => X"00000000",
		16#04c9# => X"00000000",
		16#04ca# => X"00000000",
		16#04cb# => X"00000000",
		16#04cc# => X"00000000",
		16#04cd# => X"00000000",
		16#04ce# => X"00000000",
		16#04cf# => X"00000000",
		16#04d0# => X"00000000",
		16#04d1# => X"00000000",
		16#04d2# => X"00000000",
		16#04d3# => X"00000000",
		16#04d4# => X"00000000",
		16#04d5# => X"00000000",
		16#04d6# => X"00000000",
		16#04d7# => X"00000000",
		16#04d8# => X"00000000",
		16#04d9# => X"00000000",
		16#04da# => X"00000000",
		16#04db# => X"00000000",
		16#04dc# => X"00000000",
		16#04dd# => X"00000000",
		16#04de# => X"00000000",
		16#04df# => X"00000000",
		16#04e0# => X"00000000",
		16#04e1# => X"00000000",
		16#04e2# => X"00000000",
		16#04e3# => X"00000000",
		16#04e4# => X"00000000",
		16#04e5# => X"00000000",
		16#04e6# => X"00000000",
		16#04e7# => X"00000000",
		16#04e8# => X"00000000",
		16#04e9# => X"00000000",
		16#04ea# => X"00000000",
		16#04eb# => X"00000000",
		16#04ec# => X"00000000",
		16#04ed# => X"00000000",
		16#04ee# => X"00000000",
		16#04ef# => X"00000000",
		16#04f0# => X"00000000",
		16#04f1# => X"00000000",
		16#04f2# => X"00000000",
		16#04f3# => X"00000000",
		16#04f4# => X"00000000",
		16#04f5# => X"00000000",
		16#04f6# => X"00000000",
		16#04f7# => X"00000000",
		16#04f8# => X"00000000",
		16#04f9# => X"00000000",
		16#04fa# => X"00000000",
		16#04fb# => X"00000000",
		16#04fc# => X"00000000",
		16#04fd# => X"00000000",
		16#04fe# => X"00000000",
		16#04ff# => X"00000000",
		16#0500# => X"9c21ff00",
		16#0501# => X"d4011804",
		16#0502# => X"d4012008",
		16#0503# => X"b4600010",
		16#0504# => X"00002fa4",
		16#0505# => X"b4800020",
		16#0506# => X"00000000",
		16#0507# => X"00000000",
		16#0508# => X"00000000",
		16#0509# => X"00000000",
		16#050a# => X"00000000",
		16#050b# => X"00000000",
		16#050c# => X"00000000",
		16#050d# => X"00000000",
		16#050e# => X"00000000",
		16#050f# => X"00000000",
		16#0510# => X"00000000",
		16#0511# => X"00000000",
		16#0512# => X"00000000",
		16#0513# => X"00000000",
		16#0514# => X"00000000",
		16#0515# => X"00000000",
		16#0516# => X"00000000",
		16#0517# => X"00000000",
		16#0518# => X"00000000",
		16#0519# => X"00000000",
		16#051a# => X"00000000",
		16#051b# => X"00000000",
		16#051c# => X"00000000",
		16#051d# => X"00000000",
		16#051e# => X"00000000",
		16#051f# => X"00000000",
		16#0520# => X"00000000",
		16#0521# => X"00000000",
		16#0522# => X"00000000",
		16#0523# => X"00000000",
		16#0524# => X"00000000",
		16#0525# => X"00000000",
		16#0526# => X"00000000",
		16#0527# => X"00000000",
		16#0528# => X"00000000",
		16#0529# => X"00000000",
		16#052a# => X"00000000",
		16#052b# => X"00000000",
		16#052c# => X"00000000",
		16#052d# => X"00000000",
		16#052e# => X"00000000",
		16#052f# => X"00000000",
		16#0530# => X"00000000",
		16#0531# => X"00000000",
		16#0532# => X"00000000",
		16#0533# => X"00000000",
		16#0534# => X"00000000",
		16#0535# => X"00000000",
		16#0536# => X"00000000",
		16#0537# => X"00000000",
		16#0538# => X"00000000",
		16#0539# => X"00000000",
		16#053a# => X"00000000",
		16#053b# => X"00000000",
		16#053c# => X"00000000",
		16#053d# => X"00000000",
		16#053e# => X"00000000",
		16#053f# => X"00000000",
		16#0540# => X"9c21ff00",
		16#0541# => X"d4011804",
		16#0542# => X"d4012008",
		16#0543# => X"b4600010",
		16#0544# => X"00002f64",
		16#0545# => X"b4800020",
		16#0546# => X"00000000",
		16#0547# => X"00000000",
		16#0548# => X"00000000",
		16#0549# => X"00000000",
		16#054a# => X"00000000",
		16#054b# => X"00000000",
		16#054c# => X"00000000",
		16#054d# => X"00000000",
		16#054e# => X"00000000",
		16#054f# => X"00000000",
		16#0550# => X"00000000",
		16#0551# => X"00000000",
		16#0552# => X"00000000",
		16#0553# => X"00000000",
		16#0554# => X"00000000",
		16#0555# => X"00000000",
		16#0556# => X"00000000",
		16#0557# => X"00000000",
		16#0558# => X"00000000",
		16#0559# => X"00000000",
		16#055a# => X"00000000",
		16#055b# => X"00000000",
		16#055c# => X"00000000",
		16#055d# => X"00000000",
		16#055e# => X"00000000",
		16#055f# => X"00000000",
		16#0560# => X"00000000",
		16#0561# => X"00000000",
		16#0562# => X"00000000",
		16#0563# => X"00000000",
		16#0564# => X"00000000",
		16#0565# => X"00000000",
		16#0566# => X"00000000",
		16#0567# => X"00000000",
		16#0568# => X"00000000",
		16#0569# => X"00000000",
		16#056a# => X"00000000",
		16#056b# => X"00000000",
		16#056c# => X"00000000",
		16#056d# => X"00000000",
		16#056e# => X"00000000",
		16#056f# => X"00000000",
		16#0570# => X"00000000",
		16#0571# => X"00000000",
		16#0572# => X"00000000",
		16#0573# => X"00000000",
		16#0574# => X"00000000",
		16#0575# => X"00000000",
		16#0576# => X"00000000",
		16#0577# => X"00000000",
		16#0578# => X"00000000",
		16#0579# => X"00000000",
		16#057a# => X"00000000",
		16#057b# => X"00000000",
		16#057c# => X"00000000",
		16#057d# => X"00000000",
		16#057e# => X"00000000",
		16#057f# => X"00000000",
		16#0580# => X"9c21ff00",
		16#0581# => X"d4011804",
		16#0582# => X"d4012008",
		16#0583# => X"b4600010",
		16#0584# => X"00002f24",
		16#0585# => X"b4800020",
		16#0586# => X"00000000",
		16#0587# => X"00000000",
		16#0588# => X"00000000",
		16#0589# => X"00000000",
		16#058a# => X"00000000",
		16#058b# => X"00000000",
		16#058c# => X"00000000",
		16#058d# => X"00000000",
		16#058e# => X"00000000",
		16#058f# => X"00000000",
		16#0590# => X"00000000",
		16#0591# => X"00000000",
		16#0592# => X"00000000",
		16#0593# => X"00000000",
		16#0594# => X"00000000",
		16#0595# => X"00000000",
		16#0596# => X"00000000",
		16#0597# => X"00000000",
		16#0598# => X"00000000",
		16#0599# => X"00000000",
		16#059a# => X"00000000",
		16#059b# => X"00000000",
		16#059c# => X"00000000",
		16#059d# => X"00000000",
		16#059e# => X"00000000",
		16#059f# => X"00000000",
		16#05a0# => X"00000000",
		16#05a1# => X"00000000",
		16#05a2# => X"00000000",
		16#05a3# => X"00000000",
		16#05a4# => X"00000000",
		16#05a5# => X"00000000",
		16#05a6# => X"00000000",
		16#05a7# => X"00000000",
		16#05a8# => X"00000000",
		16#05a9# => X"00000000",
		16#05aa# => X"00000000",
		16#05ab# => X"00000000",
		16#05ac# => X"00000000",
		16#05ad# => X"00000000",
		16#05ae# => X"00000000",
		16#05af# => X"00000000",
		16#05b0# => X"00000000",
		16#05b1# => X"00000000",
		16#05b2# => X"00000000",
		16#05b3# => X"00000000",
		16#05b4# => X"00000000",
		16#05b5# => X"00000000",
		16#05b6# => X"00000000",
		16#05b7# => X"00000000",
		16#05b8# => X"00000000",
		16#05b9# => X"00000000",
		16#05ba# => X"00000000",
		16#05bb# => X"00000000",
		16#05bc# => X"00000000",
		16#05bd# => X"00000000",
		16#05be# => X"00000000",
		16#05bf# => X"00000000",
		16#05c0# => X"9c21ff00",
		16#05c1# => X"d4011804",
		16#05c2# => X"d4012008",
		16#05c3# => X"b4600010",
		16#05c4# => X"00002ee4",
		16#05c5# => X"b4800020",
		16#05c6# => X"00000000",
		16#05c7# => X"00000000",
		16#05c8# => X"00000000",
		16#05c9# => X"00000000",
		16#05ca# => X"00000000",
		16#05cb# => X"00000000",
		16#05cc# => X"00000000",
		16#05cd# => X"00000000",
		16#05ce# => X"00000000",
		16#05cf# => X"00000000",
		16#05d0# => X"00000000",
		16#05d1# => X"00000000",
		16#05d2# => X"00000000",
		16#05d3# => X"00000000",
		16#05d4# => X"00000000",
		16#05d5# => X"00000000",
		16#05d6# => X"00000000",
		16#05d7# => X"00000000",
		16#05d8# => X"00000000",
		16#05d9# => X"00000000",
		16#05da# => X"00000000",
		16#05db# => X"00000000",
		16#05dc# => X"00000000",
		16#05dd# => X"00000000",
		16#05de# => X"00000000",
		16#05df# => X"00000000",
		16#05e0# => X"00000000",
		16#05e1# => X"00000000",
		16#05e2# => X"00000000",
		16#05e3# => X"00000000",
		16#05e4# => X"00000000",
		16#05e5# => X"00000000",
		16#05e6# => X"00000000",
		16#05e7# => X"00000000",
		16#05e8# => X"00000000",
		16#05e9# => X"00000000",
		16#05ea# => X"00000000",
		16#05eb# => X"00000000",
		16#05ec# => X"00000000",
		16#05ed# => X"00000000",
		16#05ee# => X"00000000",
		16#05ef# => X"00000000",
		16#05f0# => X"00000000",
		16#05f1# => X"00000000",
		16#05f2# => X"00000000",
		16#05f3# => X"00000000",
		16#05f4# => X"00000000",
		16#05f5# => X"00000000",
		16#05f6# => X"00000000",
		16#05f7# => X"00000000",
		16#05f8# => X"00000000",
		16#05f9# => X"00000000",
		16#05fa# => X"00000000",
		16#05fb# => X"00000000",
		16#05fc# => X"00000000",
		16#05fd# => X"00000000",
		16#05fe# => X"00000000",
		16#05ff# => X"00000000",
		16#0600# => X"9c21ff00",
		16#0601# => X"d4011804",
		16#0602# => X"d4012008",
		16#0603# => X"b4600010",
		16#0604# => X"00002ea4",
		16#0605# => X"b4800020",
		16#0606# => X"00000000",
		16#0607# => X"00000000",
		16#0608# => X"00000000",
		16#0609# => X"00000000",
		16#060a# => X"00000000",
		16#060b# => X"00000000",
		16#060c# => X"00000000",
		16#060d# => X"00000000",
		16#060e# => X"00000000",
		16#060f# => X"00000000",
		16#0610# => X"00000000",
		16#0611# => X"00000000",
		16#0612# => X"00000000",
		16#0613# => X"00000000",
		16#0614# => X"00000000",
		16#0615# => X"00000000",
		16#0616# => X"00000000",
		16#0617# => X"00000000",
		16#0618# => X"00000000",
		16#0619# => X"00000000",
		16#061a# => X"00000000",
		16#061b# => X"00000000",
		16#061c# => X"00000000",
		16#061d# => X"00000000",
		16#061e# => X"00000000",
		16#061f# => X"00000000",
		16#0620# => X"00000000",
		16#0621# => X"00000000",
		16#0622# => X"00000000",
		16#0623# => X"00000000",
		16#0624# => X"00000000",
		16#0625# => X"00000000",
		16#0626# => X"00000000",
		16#0627# => X"00000000",
		16#0628# => X"00000000",
		16#0629# => X"00000000",
		16#062a# => X"00000000",
		16#062b# => X"00000000",
		16#062c# => X"00000000",
		16#062d# => X"00000000",
		16#062e# => X"00000000",
		16#062f# => X"00000000",
		16#0630# => X"00000000",
		16#0631# => X"00000000",
		16#0632# => X"00000000",
		16#0633# => X"00000000",
		16#0634# => X"00000000",
		16#0635# => X"00000000",
		16#0636# => X"00000000",
		16#0637# => X"00000000",
		16#0638# => X"00000000",
		16#0639# => X"00000000",
		16#063a# => X"00000000",
		16#063b# => X"00000000",
		16#063c# => X"00000000",
		16#063d# => X"00000000",
		16#063e# => X"00000000",
		16#063f# => X"00000000",
		16#0640# => X"9c21ff00",
		16#0641# => X"d4011804",
		16#0642# => X"d4012008",
		16#0643# => X"b4600010",
		16#0644# => X"00002e64",
		16#0645# => X"b4800020",
		16#0646# => X"00000000",
		16#0647# => X"00000000",
		16#0648# => X"00000000",
		16#0649# => X"00000000",
		16#064a# => X"00000000",
		16#064b# => X"00000000",
		16#064c# => X"00000000",
		16#064d# => X"00000000",
		16#064e# => X"00000000",
		16#064f# => X"00000000",
		16#0650# => X"00000000",
		16#0651# => X"00000000",
		16#0652# => X"00000000",
		16#0653# => X"00000000",
		16#0654# => X"00000000",
		16#0655# => X"00000000",
		16#0656# => X"00000000",
		16#0657# => X"00000000",
		16#0658# => X"00000000",
		16#0659# => X"00000000",
		16#065a# => X"00000000",
		16#065b# => X"00000000",
		16#065c# => X"00000000",
		16#065d# => X"00000000",
		16#065e# => X"00000000",
		16#065f# => X"00000000",
		16#0660# => X"00000000",
		16#0661# => X"00000000",
		16#0662# => X"00000000",
		16#0663# => X"00000000",
		16#0664# => X"00000000",
		16#0665# => X"00000000",
		16#0666# => X"00000000",
		16#0667# => X"00000000",
		16#0668# => X"00000000",
		16#0669# => X"00000000",
		16#066a# => X"00000000",
		16#066b# => X"00000000",
		16#066c# => X"00000000",
		16#066d# => X"00000000",
		16#066e# => X"00000000",
		16#066f# => X"00000000",
		16#0670# => X"00000000",
		16#0671# => X"00000000",
		16#0672# => X"00000000",
		16#0673# => X"00000000",
		16#0674# => X"00000000",
		16#0675# => X"00000000",
		16#0676# => X"00000000",
		16#0677# => X"00000000",
		16#0678# => X"00000000",
		16#0679# => X"00000000",
		16#067a# => X"00000000",
		16#067b# => X"00000000",
		16#067c# => X"00000000",
		16#067d# => X"00000000",
		16#067e# => X"00000000",
		16#067f# => X"00000000",
		16#0680# => X"9c21ff00",
		16#0681# => X"d4011804",
		16#0682# => X"d4012008",
		16#0683# => X"b4600010",
		16#0684# => X"00002e24",
		16#0685# => X"b4800020",
		16#0686# => X"00000000",
		16#0687# => X"00000000",
		16#0688# => X"00000000",
		16#0689# => X"00000000",
		16#068a# => X"00000000",
		16#068b# => X"00000000",
		16#068c# => X"00000000",
		16#068d# => X"00000000",
		16#068e# => X"00000000",
		16#068f# => X"00000000",
		16#0690# => X"00000000",
		16#0691# => X"00000000",
		16#0692# => X"00000000",
		16#0693# => X"00000000",
		16#0694# => X"00000000",
		16#0695# => X"00000000",
		16#0696# => X"00000000",
		16#0697# => X"00000000",
		16#0698# => X"00000000",
		16#0699# => X"00000000",
		16#069a# => X"00000000",
		16#069b# => X"00000000",
		16#069c# => X"00000000",
		16#069d# => X"00000000",
		16#069e# => X"00000000",
		16#069f# => X"00000000",
		16#06a0# => X"00000000",
		16#06a1# => X"00000000",
		16#06a2# => X"00000000",
		16#06a3# => X"00000000",
		16#06a4# => X"00000000",
		16#06a5# => X"00000000",
		16#06a6# => X"00000000",
		16#06a7# => X"00000000",
		16#06a8# => X"00000000",
		16#06a9# => X"00000000",
		16#06aa# => X"00000000",
		16#06ab# => X"00000000",
		16#06ac# => X"00000000",
		16#06ad# => X"00000000",
		16#06ae# => X"00000000",
		16#06af# => X"00000000",
		16#06b0# => X"00000000",
		16#06b1# => X"00000000",
		16#06b2# => X"00000000",
		16#06b3# => X"00000000",
		16#06b4# => X"00000000",
		16#06b5# => X"00000000",
		16#06b6# => X"00000000",
		16#06b7# => X"00000000",
		16#06b8# => X"00000000",
		16#06b9# => X"00000000",
		16#06ba# => X"00000000",
		16#06bb# => X"00000000",
		16#06bc# => X"00000000",
		16#06bd# => X"00000000",
		16#06be# => X"00000000",
		16#06bf# => X"00000000",
		16#06c0# => X"9c21ff00",
		16#06c1# => X"d4011804",
		16#06c2# => X"d4012008",
		16#06c3# => X"b4600010",
		16#06c4# => X"00002de4",
		16#06c5# => X"b4800020",
		16#06c6# => X"00000000",
		16#06c7# => X"00000000",
		16#06c8# => X"00000000",
		16#06c9# => X"00000000",
		16#06ca# => X"00000000",
		16#06cb# => X"00000000",
		16#06cc# => X"00000000",
		16#06cd# => X"00000000",
		16#06ce# => X"00000000",
		16#06cf# => X"00000000",
		16#06d0# => X"00000000",
		16#06d1# => X"00000000",
		16#06d2# => X"00000000",
		16#06d3# => X"00000000",
		16#06d4# => X"00000000",
		16#06d5# => X"00000000",
		16#06d6# => X"00000000",
		16#06d7# => X"00000000",
		16#06d8# => X"00000000",
		16#06d9# => X"00000000",
		16#06da# => X"00000000",
		16#06db# => X"00000000",
		16#06dc# => X"00000000",
		16#06dd# => X"00000000",
		16#06de# => X"00000000",
		16#06df# => X"00000000",
		16#06e0# => X"00000000",
		16#06e1# => X"00000000",
		16#06e2# => X"00000000",
		16#06e3# => X"00000000",
		16#06e4# => X"00000000",
		16#06e5# => X"00000000",
		16#06e6# => X"00000000",
		16#06e7# => X"00000000",
		16#06e8# => X"00000000",
		16#06e9# => X"00000000",
		16#06ea# => X"00000000",
		16#06eb# => X"00000000",
		16#06ec# => X"00000000",
		16#06ed# => X"00000000",
		16#06ee# => X"00000000",
		16#06ef# => X"00000000",
		16#06f0# => X"00000000",
		16#06f1# => X"00000000",
		16#06f2# => X"00000000",
		16#06f3# => X"00000000",
		16#06f4# => X"00000000",
		16#06f5# => X"00000000",
		16#06f6# => X"00000000",
		16#06f7# => X"00000000",
		16#06f8# => X"00000000",
		16#06f9# => X"00000000",
		16#06fa# => X"00000000",
		16#06fb# => X"00000000",
		16#06fc# => X"00000000",
		16#06fd# => X"00000000",
		16#06fe# => X"00000000",
		16#06ff# => X"00000000",
		16#0700# => X"9c21ff00",
		16#0701# => X"d4011804",
		16#0702# => X"d4012008",
		16#0703# => X"b4600010",
		16#0704# => X"00002da4",
		16#0705# => X"b4800020",
		16#0706# => X"00000000",
		16#0707# => X"00000000",
		16#0708# => X"00000000",
		16#0709# => X"00000000",
		16#070a# => X"00000000",
		16#070b# => X"00000000",
		16#070c# => X"00000000",
		16#070d# => X"00000000",
		16#070e# => X"00000000",
		16#070f# => X"00000000",
		16#0710# => X"00000000",
		16#0711# => X"00000000",
		16#0712# => X"00000000",
		16#0713# => X"00000000",
		16#0714# => X"00000000",
		16#0715# => X"00000000",
		16#0716# => X"00000000",
		16#0717# => X"00000000",
		16#0718# => X"00000000",
		16#0719# => X"00000000",
		16#071a# => X"00000000",
		16#071b# => X"00000000",
		16#071c# => X"00000000",
		16#071d# => X"00000000",
		16#071e# => X"00000000",
		16#071f# => X"00000000",
		16#0720# => X"00000000",
		16#0721# => X"00000000",
		16#0722# => X"00000000",
		16#0723# => X"00000000",
		16#0724# => X"00000000",
		16#0725# => X"00000000",
		16#0726# => X"00000000",
		16#0727# => X"00000000",
		16#0728# => X"00000000",
		16#0729# => X"00000000",
		16#072a# => X"00000000",
		16#072b# => X"00000000",
		16#072c# => X"00000000",
		16#072d# => X"00000000",
		16#072e# => X"00000000",
		16#072f# => X"00000000",
		16#0730# => X"00000000",
		16#0731# => X"00000000",
		16#0732# => X"00000000",
		16#0733# => X"00000000",
		16#0734# => X"00000000",
		16#0735# => X"00000000",
		16#0736# => X"00000000",
		16#0737# => X"00000000",
		16#0738# => X"00000000",
		16#0739# => X"00000000",
		16#073a# => X"00000000",
		16#073b# => X"00000000",
		16#073c# => X"00000000",
		16#073d# => X"00000000",
		16#073e# => X"00000000",
		16#073f# => X"00000000",
		16#0740# => X"9c21ff00",
		16#0741# => X"d4011804",
		16#0742# => X"d4012008",
		16#0743# => X"b4600010",
		16#0744# => X"00002d64",
		16#0745# => X"b4800020",
		16#0746# => X"00000000",
		16#0747# => X"00000000",
		16#0748# => X"00000000",
		16#0749# => X"00000000",
		16#074a# => X"00000000",
		16#074b# => X"00000000",
		16#074c# => X"00000000",
		16#074d# => X"00000000",
		16#074e# => X"00000000",
		16#074f# => X"00000000",
		16#0750# => X"00000000",
		16#0751# => X"00000000",
		16#0752# => X"00000000",
		16#0753# => X"00000000",
		16#0754# => X"00000000",
		16#0755# => X"00000000",
		16#0756# => X"00000000",
		16#0757# => X"00000000",
		16#0758# => X"00000000",
		16#0759# => X"00000000",
		16#075a# => X"00000000",
		16#075b# => X"00000000",
		16#075c# => X"00000000",
		16#075d# => X"00000000",
		16#075e# => X"00000000",
		16#075f# => X"00000000",
		16#0760# => X"00000000",
		16#0761# => X"00000000",
		16#0762# => X"00000000",
		16#0763# => X"00000000",
		16#0764# => X"00000000",
		16#0765# => X"00000000",
		16#0766# => X"00000000",
		16#0767# => X"00000000",
		16#0768# => X"00000000",
		16#0769# => X"00000000",
		16#076a# => X"00000000",
		16#076b# => X"00000000",
		16#076c# => X"00000000",
		16#076d# => X"00000000",
		16#076e# => X"00000000",
		16#076f# => X"00000000",
		16#0770# => X"00000000",
		16#0771# => X"00000000",
		16#0772# => X"00000000",
		16#0773# => X"00000000",
		16#0774# => X"00000000",
		16#0775# => X"00000000",
		16#0776# => X"00000000",
		16#0777# => X"00000000",
		16#0778# => X"00000000",
		16#0779# => X"00000000",
		16#077a# => X"00000000",
		16#077b# => X"00000000",
		16#077c# => X"00000000",
		16#077d# => X"00000000",
		16#077e# => X"00000000",
		16#077f# => X"00000000",
		16#0780# => X"9c21ff00",
		16#0781# => X"d4011804",
		16#0782# => X"d4012008",
		16#0783# => X"b4600010",
		16#0784# => X"00002d24",
		16#0785# => X"b4800020",
		16#0786# => X"00000000",
		16#0787# => X"00000000",
		16#0788# => X"00000000",
		16#0789# => X"00000000",
		16#078a# => X"00000000",
		16#078b# => X"00000000",
		16#078c# => X"00000000",
		16#078d# => X"00000000",
		16#078e# => X"00000000",
		16#078f# => X"00000000",
		16#0790# => X"00000000",
		16#0791# => X"00000000",
		16#0792# => X"00000000",
		16#0793# => X"00000000",
		16#0794# => X"00000000",
		16#0795# => X"00000000",
		16#0796# => X"00000000",
		16#0797# => X"00000000",
		16#0798# => X"00000000",
		16#0799# => X"00000000",
		16#079a# => X"00000000",
		16#079b# => X"00000000",
		16#079c# => X"00000000",
		16#079d# => X"00000000",
		16#079e# => X"00000000",
		16#079f# => X"00000000",
		16#07a0# => X"00000000",
		16#07a1# => X"00000000",
		16#07a2# => X"00000000",
		16#07a3# => X"00000000",
		16#07a4# => X"00000000",
		16#07a5# => X"00000000",
		16#07a6# => X"00000000",
		16#07a7# => X"00000000",
		16#07a8# => X"00000000",
		16#07a9# => X"00000000",
		16#07aa# => X"00000000",
		16#07ab# => X"00000000",
		16#07ac# => X"00000000",
		16#07ad# => X"00000000",
		16#07ae# => X"00000000",
		16#07af# => X"00000000",
		16#07b0# => X"00000000",
		16#07b1# => X"00000000",
		16#07b2# => X"00000000",
		16#07b3# => X"00000000",
		16#07b4# => X"00000000",
		16#07b5# => X"00000000",
		16#07b6# => X"00000000",
		16#07b7# => X"00000000",
		16#07b8# => X"00000000",
		16#07b9# => X"00000000",
		16#07ba# => X"00000000",
		16#07bb# => X"00000000",
		16#07bc# => X"00000000",
		16#07bd# => X"00000000",
		16#07be# => X"00000000",
		16#07bf# => X"00000000",
		16#07c0# => X"9c21ff00",
		16#07c1# => X"d4011804",
		16#07c2# => X"d4012008",
		16#07c3# => X"b4600010",
		16#07c4# => X"00002ce4",
		16#07c5# => X"b4800020",
		16#07c6# => X"00000000",
		16#07c7# => X"00000000",
		16#07c8# => X"00000000",
		16#07c9# => X"00000000",
		16#07ca# => X"00000000",
		16#07cb# => X"00000000",
		16#07cc# => X"00000000",
		16#07cd# => X"00000000",
		16#07ce# => X"00000000",
		16#07cf# => X"00000000",
		16#07d0# => X"00000000",
		16#07d1# => X"00000000",
		16#07d2# => X"00000000",
		16#07d3# => X"00000000",
		16#07d4# => X"00000000",
		16#07d5# => X"00000000",
		16#07d6# => X"00000000",
		16#07d7# => X"00000000",
		16#07d8# => X"00000000",
		16#07d9# => X"00000000",
		16#07da# => X"00000000",
		16#07db# => X"00000000",
		16#07dc# => X"00000000",
		16#07dd# => X"00000000",
		16#07de# => X"00000000",
		16#07df# => X"00000000",
		16#07e0# => X"00000000",
		16#07e1# => X"00000000",
		16#07e2# => X"00000000",
		16#07e3# => X"00000000",
		16#07e4# => X"00000000",
		16#07e5# => X"00000000",
		16#07e6# => X"00000000",
		16#07e7# => X"00000000",
		16#07e8# => X"00000000",
		16#07e9# => X"00000000",
		16#07ea# => X"00000000",
		16#07eb# => X"00000000",
		16#07ec# => X"00000000",
		16#07ed# => X"00000000",
		16#07ee# => X"00000000",
		16#07ef# => X"00000000",
		16#07f0# => X"00000000",
		16#07f1# => X"00000000",
		16#07f2# => X"00000000",
		16#07f3# => X"00000000",
		16#07f4# => X"00000000",
		16#07f5# => X"00000000",
		16#07f6# => X"00000000",
		16#07f7# => X"00000000",
		16#07f8# => X"00000000",
		16#07f9# => X"00000000",
		16#07fa# => X"00000000",
		16#07fb# => X"00000000",
		16#07fc# => X"00000000",
		16#07fd# => X"00000000",
		16#07fe# => X"00000000",
		16#07ff# => X"15000000",
		16#0800# => X"15000000",
		16#0801# => X"9c21fffc",
		16#0802# => X"d4014800",
		16#0803# => X"04000071",
		16#0804# => X"15000000",
		16#0805# => X"0400578a",
		16#0806# => X"15000000",
		16#0807# => X"85210000",
		16#0808# => X"44004800",
		16#0809# => X"9c210004",
		16#080a# => X"18200001",
		16#080b# => X"a8217d9c",
		16#080c# => X"84210000",
		16#080d# => X"18400001",
		16#080e# => X"a8427da0",
		16#080f# => X"84420000",
		16#0810# => X"e0211000",
		16#0811# => X"e0410804",
		16#0812# => X"b460c002",
		16#0813# => X"b0838000",
		16#0814# => X"e0212000",
		16#0815# => X"18600001",
		16#0816# => X"a863adc4",
		16#0817# => X"d4030800",
		16#0818# => X"04002be2",
		16#0819# => X"15000000",
		16#081a# => X"18600001",
		16#081b# => X"a863b7e0",
		16#081c# => X"18800001",
		16#081d# => X"a884c50c",
		16#081e# => X"d4030000",
		16#081f# => X"e4832000",
		16#0820# => X"13fffffe",
		16#0821# => X"9c630004",
		16#0822# => X"040055c6",
		16#0823# => X"15000000",
		16#0824# => X"07ffffdd",
		16#0825# => X"15000000",
		16#0826# => X"18600001",
		16#0827# => X"04002935",
		16#0828# => X"a8637ea0",
		16#0829# => X"18800001",
		16#082a# => X"a8847da8",
		16#082b# => X"84840000",
		16#082c# => X"e4240000",
		16#082d# => X"0c000004",
		16#082e# => X"e0600004",
		16#082f# => X"040056b1",
		16#0830# => X"15000000",
		16#0831# => X"e0600004",
		16#0832# => X"e0800004",
		16#0833# => X"0400044d",
		16#0834# => X"e0a00004",
		16#0835# => X"04002930",
		16#0836# => X"9c6b0000",
		16#0837# => X"00000000",
		16#0838# => X"15000000",
		16#0839# => X"d7e187f8",
		16#083a# => X"1a000001",
		16#083b# => X"d7e117f0",
		16#083c# => X"aa10b7e0",
		16#083d# => X"d7e14ffc",
		16#083e# => X"8c500000",
		16#083f# => X"d7e177f4",
		16#0840# => X"bc220000",
		16#0841# => X"10000027",
		16#0842# => X"9c21fff0",
		16#0843# => X"19c00001",
		16#0844# => X"18800001",
		16#0845# => X"a9ceadbc",
		16#0846# => X"a884adb8",
		16#0847# => X"18400001",
		16#0848# => X"e1ce2002",
		16#0849# => X"a842b7e4",
		16#084a# => X"b9ce0082",
		16#084b# => X"84620000",
		16#084c# => X"9dceffff",
		16#084d# => X"e4637000",
		16#084e# => X"10000010",
		16#084f# => X"15000000",
		16#0850# => X"9c630001",
		16#0851# => X"18a00001",
		16#0852# => X"b8830002",
		16#0853# => X"a8a5adb8",
		16#0854# => X"d4021800",
		16#0855# => X"e0642800",
		16#0856# => X"84630000",
		16#0857# => X"48001800",
		16#0858# => X"15000000",
		16#0859# => X"84620000",
		16#085a# => X"e4837000",
		16#085b# => X"13fffff6",
		16#085c# => X"9c630001",
		16#085d# => X"9c63ffff",
		16#085e# => X"18400000",
		16#085f# => X"a8420000",
		16#0860# => X"bc020000",
		16#0861# => X"10000006",
		16#0862# => X"9c400001",
		16#0863# => X"18600001",
		16#0864# => X"07fff79c",
		16#0865# => X"a8638dac",
		16#0866# => X"9c400001",
		16#0867# => X"d8101000",
		16#0868# => X"9c210010",
		16#0869# => X"8521fffc",
		16#086a# => X"8441fff0",
		16#086b# => X"85c1fff4",
		16#086c# => X"44004800",
		16#086d# => X"8601fff8",
		16#086e# => X"d7e14ffc",
		16#086f# => X"9c21fffc",
		16#0870# => X"9c210004",
		16#0871# => X"8521fffc",
		16#0872# => X"44004800",
		16#0873# => X"15000000",
		16#0874# => X"18600000",
		16#0875# => X"d7e14ffc",
		16#0876# => X"a8630000",
		16#0877# => X"bc030000",
		16#0878# => X"10000007",
		16#0879# => X"9c21fffc",
		16#087a# => X"18600001",
		16#087b# => X"18800001",
		16#087c# => X"a8638dac",
		16#087d# => X"07fff783",
		16#087e# => X"a884b7e8",
		16#087f# => X"18600001",
		16#0880# => X"a863adc0",
		16#0881# => X"84830000",
		16#0882# => X"bc040000",
		16#0883# => X"1000000a",
		16#0884# => X"18800000",
		16#0885# => X"a8840000",
		16#0886# => X"bc040000",
		16#0887# => X"10000006",
		16#0888# => X"15000000",
		16#0889# => X"9c210004",
		16#088a# => X"8521fffc",
		16#088b# => X"44002000",
		16#088c# => X"15000000",
		16#088d# => X"9c210004",
		16#088e# => X"8521fffc",
		16#088f# => X"44004800",
		16#0890# => X"15000000",
		16#0891# => X"d7e14ffc",
		16#0892# => X"9c21fffc",
		16#0893# => X"9c210004",
		16#0894# => X"8521fffc",
		16#0895# => X"44004800",
		16#0896# => X"15000000",
		16#0897# => X"d7e117fc",
		16#0898# => X"bc250000",
		16#0899# => X"0c000008",
		16#089a# => X"9c21fffc",
		16#089b# => X"99630002",
		16#089c# => X"98640002",
		16#089d# => X"9c210004",
		16#089e# => X"e16b1802",
		16#089f# => X"44004800",
		16#08a0# => X"8441fffc",
		16#08a1# => X"98a30000",
		16#08a2# => X"a4c5ffff",
		16#08a3# => X"9c40ff00",
		16#08a4# => X"b8c60048",
		16#08a5# => X"e0a51003",
		16#08a6# => X"99630002",
		16#08a7# => X"e0a62804",
		16#08a8# => X"dc032800",
		16#08a9# => X"98640002",
		16#08aa# => X"98a40000",
		16#08ab# => X"a4c5ffff",
		16#08ac# => X"e0a51003",
		16#08ad# => X"b8c60048",
		16#08ae# => X"9c210004",
		16#08af# => X"e16b1802",
		16#08b0# => X"e0a62804",
		16#08b1# => X"8441fffc",
		16#08b2# => X"44004800",
		16#08b3# => X"dc042800",
		16#08b4# => X"d7e177f0",
		16#08b5# => X"99c30000",
		16#08b6# => X"d7e197f8",
		16#08b7# => X"aa430000",
		16#08b8# => X"b86e0087",
		16#08b9# => X"d7e117ec",
		16#08ba# => X"d7e14ffc",
		16#08bb# => X"d7e187f4",
		16#08bc# => X"a4630001",
		16#08bd# => X"9c21ffec",
		16#08be# => X"bc030000",
		16#08bf# => X"0c00002e",
		16#08c0# => X"a8440000",
		16#08c1# => X"b88e0043",
		16#08c2# => X"a46e0007",
		16#08c3# => X"a484000f",
		16#08c4# => X"bc030000",
		16#08c5# => X"b8a40004",
		16#08c6# => X"10000017",
		16#08c7# => X"e0852004",
		16#08c8# => X"bc030001",
		16#08c9# => X"1000002d",
		16#08ca# => X"aa0e0000",
		16#08cb# => X"94820038",
		16#08cc# => X"04000fef",
		16#08cd# => X"a470ffff",
		16#08ce# => X"9c60ff00",
		16#08cf# => X"a490007f",
		16#08d0# => X"e1ce1803",
		16#08d1# => X"dc025838",
		16#08d2# => X"a9ce0080",
		16#08d3# => X"a9640000",
		16#08d4# => X"e1c47004",
		16#08d5# => X"dc127000",
		16#08d6# => X"9c210014",
		16#08d7# => X"8521fffc",
		16#08d8# => X"8441ffec",
		16#08d9# => X"85c1fff0",
		16#08da# => X"8601fff4",
		16#08db# => X"44004800",
		16#08dc# => X"8641fff8",
		16#08dd# => X"bda40021",
		16#08de# => X"0c000022",
		16#08df# => X"9ce00022",
		16#08e0# => X"98a20000",
		16#08e1# => X"98c20002",
		16#08e2# => X"95020038",
		16#08e3# => X"84620018",
		16#08e4# => X"04000ea6",
		16#08e5# => X"84820014",
		16#08e6# => X"9462003e",
		16#08e7# => X"ba0b0010",
		16#08e8# => X"bc230000",
		16#08e9# => X"13ffffe2",
		16#08ea# => X"ba100090",
		16#08eb# => X"03ffffe0",
		16#08ec# => X"dc02583e",
		16#08ed# => X"9c210014",
		16#08ee# => X"a48e007f",
		16#08ef# => X"8521fffc",
		16#08f0# => X"a9640000",
		16#08f1# => X"8441ffec",
		16#08f2# => X"85c1fff0",
		16#08f3# => X"8601fff4",
		16#08f4# => X"44004800",
		16#08f5# => X"8641fff8",
		16#08f6# => X"94a20038",
		16#08f7# => X"04000bf2",
		16#08f8# => X"9c620028",
		16#08f9# => X"9462003c",
		16#08fa# => X"ba0b0010",
		16#08fb# => X"bc230000",
		16#08fc# => X"13ffffcf",
		16#08fd# => X"ba100090",
		16#08fe# => X"03ffffcd",
		16#08ff# => X"dc02583c",
		16#0900# => X"03ffffe0",
		16#0901# => X"a8e40000",
		16#0902# => X"d7e14ffc",
		16#0903# => X"d7e117f0",
		16#0904# => X"d7e177f4",
		16#0905# => X"d7e187f8",
		16#0906# => X"9c21fff0",
		16#0907# => X"aa040000",
		16#0908# => X"a8850000",
		16#0909# => X"07ffffab",
		16#090a# => X"a8450000",
		16#090b# => X"a8700000",
		16#090c# => X"a8820000",
		16#090d# => X"07ffffa7",
		16#090e# => X"a9cb0000",
		16#090f# => X"9c210010",
		16#0910# => X"e16e5802",
		16#0911# => X"8521fffc",
		16#0912# => X"8441fff0",
		16#0913# => X"85c1fff4",
		16#0914# => X"44004800",
		16#0915# => X"8601fff8",
		16#0916# => X"d7e117fc",
		16#0917# => X"9c21fffc",
		16#0918# => X"94440000",
		16#0919# => X"94840002",
		16#091a# => X"9c210004",
		16#091b# => X"dc031000",
		16#091c# => X"dc032002",
		16#091d# => X"44004800",
		16#091e# => X"8441fffc",
		16#091f# => X"d7e117d4",
		16#0920# => X"d7e177d8",
		16#0921# => X"d7e14ffc",
		16#0922# => X"d7e187dc",
		16#0923# => X"d7e197e0",
		16#0924# => X"d7e1a7e4",
		16#0925# => X"d7e1b7e8",
		16#0926# => X"d7e1c7ec",
		16#0927# => X"d7e1d7f0",
		16#0928# => X"d7e1e7f4",
		16#0929# => X"d7e1f7f8",
		16#092a# => X"9c21ffc0",
		16#092b# => X"b8840010",
		16#092c# => X"99a30004",
		16#092d# => X"d4011800",
		16#092e# => X"b9c40090",
		16#092f# => X"bdad0000",
		16#0930# => X"1000016d",
		16#0931# => X"84430024",
		16#0932# => X"9c600000",
		16#0933# => X"ab8e0000",
		16#0934# => X"a9830000",
		16#0935# => X"a9030000",
		16#0936# => X"a9630000",
		16#0937# => X"a48300ff",
		16#0938# => X"bd7c0000",
		16#0939# => X"0c0000bc",
		16#093a# => X"d401200c",
		16#093b# => X"bc020000",
		16#093c# => X"100000ce",
		16#093d# => X"15000000",
		16#093e# => X"84820004",
		16#093f# => X"98840002",
		16#0940# => X"e404e000",
		16#0941# => X"0c000009",
		16#0942# => X"a8a20000",
		16#0943# => X"0000000e",
		16#0944# => X"9ce00000",
		16#0945# => X"84850004",
		16#0946# => X"98c40002",
		16#0947# => X"e426e000",
		16#0948# => X"0c000009",
		16#0949# => X"15000000",
		16#094a# => X"84a50000",
		16#094b# => X"bc050000",
		16#094c# => X"0ffffff9",
		16#094d# => X"9ce00000",
		16#094e# => X"00000003",
		16#094f# => X"15000000",
		16#0950# => X"a8460000",
		16#0951# => X"84c20000",
		16#0952# => X"d4023800",
		16#0953# => X"bc260000",
		16#0954# => X"13fffffc",
		16#0955# => X"a8e20000",
		16#0956# => X"bc250000",
		16#0957# => X"0c0000b3",
		16#0958# => X"15000000",
		16#0959# => X"84850004",
		16#095a# => X"9d080001",
		16#095b# => X"98840000",
		16#095c# => X"a4c40001",
		16#095d# => X"bc060000",
		16#095e# => X"10000006",
		16#095f# => X"a508ffff",
		16#0960# => X"b8840089",
		16#0961# => X"a4840001",
		16#0962# => X"e16b2000",
		16#0963# => X"a56bffff",
		16#0964# => X"84850000",
		16#0965# => X"bc040000",
		16#0966# => X"10000008",
		16#0967# => X"bd9c0000",
		16#0968# => X"84c40000",
		16#0969# => X"d4053000",
		16#096a# => X"84a20000",
		16#096b# => X"d4042800",
		16#096c# => X"d4022000",
		16#096d# => X"bd9c0000",
		16#096e# => X"10000005",
		16#096f# => X"15000000",
		16#0970# => X"9f9c0001",
		16#0971# => X"bb9c0010",
		16#0972# => X"bb9c0090",
		16#0973# => X"9c630001",
		16#0974# => X"b8630010",
		16#0975# => X"b8630090",
		16#0976# => X"e4236800",
		16#0977# => X"13ffffc1",
		16#0978# => X"a48300ff",
		16#0979# => X"b9080002",
		16#097a# => X"bdae0000",
		16#097b# => X"e1886002",
		16#097c# => X"e16b6000",
		16#097d# => X"a56bffff",
		16#097e# => X"10000037",
		16#097f# => X"d4015810",
		16#0980# => X"bc020000",
		16#0981# => X"10000033",
		16#0982# => X"9e400001",
		16#0983# => X"9e800000",
		16#0984# => X"aa020000",
		16#0985# => X"abd40000",
		16#0986# => X"a8540000",
		16#0987# => X"9fde0001",
		16#0988# => X"a8b00000",
		16#0989# => X"9dc00000",
		16#098a# => X"84a50000",
		16#098b# => X"bc250000",
		16#098c# => X"0c000005",
		16#098d# => X"9dce0001",
		16#098e# => X"e58e9000",
		16#098f# => X"13fffffb",
		16#0990# => X"15000000",
		16#0991# => X"ab100000",
		16#0992# => X"aad20000",
		16#0993# => X"aa050000",
		16#0994# => X"bc2e0000",
		16#0995# => X"0c000011",
		16#0996# => X"e3402802",
		16#0997# => X"e0b0d004",
		16#0998# => X"bd650000",
		16#0999# => X"0c000041",
		16#099a# => X"15000000",
		16#099b# => X"a8b80000",
		16#099c# => X"9dceffff",
		16#099d# => X"87180000",
		16#099e# => X"bc140000",
		16#099f# => X"10000038",
		16#09a0# => X"15000000",
		16#09a1# => X"d4142800",
		16#09a2# => X"aa850000",
		16#09a3# => X"bc2e0000",
		16#09a4# => X"13fffff4",
		16#09a5# => X"e0b0d004",
		16#09a6# => X"e350d004",
		16#09a7# => X"bd7a0000",
		16#09a8# => X"0c000049",
		16#09a9# => X"bd560000",
		16#09aa# => X"bc300000",
		16#09ab# => X"13ffffdd",
		16#09ac# => X"9fde0001",
		16#09ad# => X"9fdeffff",
		16#09ae# => X"bc3e0001",
		16#09af# => X"0c000006",
		16#09b0# => X"d4148000",
		16#09b1# => X"bc020000",
		16#09b2# => X"0fffffd1",
		16#09b3# => X"e2529000",
		16#09b4# => X"d4021000",
		16#09b5# => X"84620000",
		16#09b6# => X"bd7c0000",
		16#09b7# => X"86030000",
		16#09b8# => X"84830004",
		16#09b9# => X"84b00000",
		16#09ba# => X"84d00004",
		16#09bb# => X"d4032800",
		16#09bc# => X"9ca00000",
		16#09bd# => X"d4033004",
		16#09be# => X"d4102004",
		16#09bf# => X"0c0000cb",
		16#09c0# => X"d4102800",
		16#09c1# => X"84620004",
		16#09c2# => X"98830002",
		16#09c3# => X"e404e000",
		16#09c4# => X"100000de",
		16#09c5# => X"15000000",
		16#09c6# => X"00000007",
		16#09c7# => X"a9c20000",
		16#09c8# => X"848e0004",
		16#09c9# => X"98840002",
		16#09ca# => X"e424e000",
		16#09cb# => X"0c000049",
		16#09cc# => X"15000000",
		16#09cd# => X"85ce0000",
		16#09ce# => X"bc0e0000",
		16#09cf# => X"0ffffff9",
		16#09d0# => X"15000000",
		16#09d1# => X"84820000",
		16#09d2# => X"bc240000",
		16#09d3# => X"10000041",
		16#09d4# => X"a9c40000",
		16#09d5# => X"00000048",
		16#09d6# => X"84c40000",
		16#09d7# => X"a8450000",
		16#09d8# => X"03ffffcb",
		16#09d9# => X"aa850000",
		16#09da# => X"e060b002",
		16#09db# => X"e063b004",
		16#09dc# => X"bd830000",
		16#09dd# => X"0fffffbf",
		16#09de# => X"a8b80000",
		16#09df# => X"84700004",
		16#09e0# => X"84810000",
		16#09e1# => X"d4011804",
		16#09e2# => X"07fffed2",
		16#09e3# => X"84780004",
		16#09e4# => X"84610004",
		16#09e5# => X"84810000",
		16#09e6# => X"07fffece",
		16#09e7# => X"d4015808",
		16#09e8# => X"84810008",
		16#09e9# => X"e0645802",
		16#09ea# => X"bd430000",
		16#09eb# => X"0fffffb0",
		16#09ec# => X"a8b00000",
		16#09ed# => X"86100000",
		16#09ee# => X"9ed6ffff",
		16#09ef# => X"03ffffaf",
		16#09f0# => X"e3408002",
		16#09f1# => X"0fffffba",
		16#09f2# => X"bc300000",
		16#09f3# => X"03fffffa",
		16#09f4# => X"a8b00000",
		16#09f5# => X"bc020000",
		16#09f6# => X"10000014",
		16#09f7# => X"84c1000c",
		16#09f8# => X"84820004",
		16#09f9# => X"8c840001",
		16#09fa# => X"e4243000",
		16#09fb# => X"10000009",
		16#09fc# => X"a8a20000",
		16#09fd# => X"03ffff54",
		16#09fe# => X"9ce00000",
		16#09ff# => X"84850004",
		16#0a00# => X"8c840001",
		16#0a01# => X"e4243000",
		16#0a02# => X"0fffff4f",
		16#0a03# => X"9ce00000",
		16#0a04# => X"84a50000",
		16#0a05# => X"bc050000",
		16#0a06# => X"0ffffff9",
		16#0a07# => X"84c1000c",
		16#0a08# => X"03ffff49",
		16#0a09# => X"9ce00000",
		16#0a0a# => X"84820000",
		16#0a0b# => X"9d8c0001",
		16#0a0c# => X"84840004",
		16#0a0d# => X"a58cffff",
		16#0a0e# => X"90840000",
		16#0a0f# => X"a4840001",
		16#0a10# => X"e16b2000",
		16#0a11# => X"03ffff5c",
		16#0a12# => X"a56bffff",
		16#0a13# => X"84620004",
		16#0a14# => X"98630000",
		16#0a15# => X"040010be",
		16#0a16# => X"84810010",
		16#0a17# => X"85ce0000",
		16#0a18# => X"bc2e0000",
		16#0a19# => X"13fffffa",
		16#0a1a# => X"d4015810",
		16#0a1b# => X"84820000",
		16#0a1c# => X"84c40000",
		16#0a1d# => X"84a40004",
		16#0a1e# => X"84700004",
		16#0a1f# => X"d4103000",
		16#0a20# => X"d4102804",
		16#0a21# => X"d4041804",
		16#0a22# => X"d4048000",
		16#0a23# => X"bc020000",
		16#0a24# => X"10000033",
		16#0a25# => X"9cc00001",
		16#0a26# => X"9e000000",
		16#0a27# => X"a8f00000",
		16#0a28# => X"a9d00000",
		16#0a29# => X"9dce0001",
		16#0a2a# => X"a8a20000",
		16#0a2b# => X"9c600000",
		16#0a2c# => X"84a50000",
		16#0a2d# => X"bc250000",
		16#0a2e# => X"0c000005",
		16#0a2f# => X"9c630001",
		16#0a30# => X"e5833000",
		16#0a31# => X"13fffffb",
		16#0a32# => X"15000000",
		16#0a33# => X"a9820000",
		16#0a34# => X"a9060000",
		16#0a35# => X"a8450000",
		16#0a36# => X"bc230000",
		16#0a37# => X"0c000011",
		16#0a38# => X"e1a02802",
		16#0a39# => X"e0a26804",
		16#0a3a# => X"bd650000",
		16#0a3b# => X"0c00002e",
		16#0a3c# => X"e0a04002",
		16#0a3d# => X"a8ac0000",
		16#0a3e# => X"9c63ffff",
		16#0a3f# => X"858c0000",
		16#0a40# => X"bc070000",
		16#0a41# => X"10000025",
		16#0a42# => X"15000000",
		16#0a43# => X"d4072800",
		16#0a44# => X"a8e50000",
		16#0a45# => X"bc230000",
		16#0a46# => X"13fffff4",
		16#0a47# => X"e0a26804",
		16#0a48# => X"e1a26804",
		16#0a49# => X"bd6d0000",
		16#0a4a# => X"0c00003c",
		16#0a4b# => X"bd480000",
		16#0a4c# => X"bc220000",
		16#0a4d# => X"13ffffdd",
		16#0a4e# => X"9dce0001",
		16#0a4f# => X"9dceffff",
		16#0a50# => X"bc2e0001",
		16#0a51# => X"0c000053",
		16#0a52# => X"d4071000",
		16#0a53# => X"a8500000",
		16#0a54# => X"bc020000",
		16#0a55# => X"0fffffd1",
		16#0a56# => X"e0c63000",
		16#0a57# => X"d4021000",
		16#0a58# => X"85610010",
		16#0a59# => X"9c210040",
		16#0a5a# => X"8521fffc",
		16#0a5b# => X"8441ffd4",
		16#0a5c# => X"85c1ffd8",
		16#0a5d# => X"8601ffdc",
		16#0a5e# => X"8641ffe0",
		16#0a5f# => X"8681ffe4",
		16#0a60# => X"86c1ffe8",
		16#0a61# => X"8701ffec",
		16#0a62# => X"8741fff0",
		16#0a63# => X"8781fff4",
		16#0a64# => X"44004800",
		16#0a65# => X"87c1fff8",
		16#0a66# => X"aa050000",
		16#0a67# => X"03ffffde",
		16#0a68# => X"a8e50000",
		16#0a69# => X"e0a54004",
		16#0a6a# => X"bd850000",
		16#0a6b# => X"0fffffd3",
		16#0a6c# => X"a8ac0000",
		16#0a6d# => X"85ec0004",
		16#0a6e# => X"9c80ff00",
		16#0a6f# => X"9a2f0000",
		16#0a70# => X"a651ffff",
		16#0a71# => X"e2312003",
		16#0a72# => X"ba520048",
		16#0a73# => X"84a20004",
		16#0a74# => X"9a6f0002",
		16#0a75# => X"e2328804",
		16#0a76# => X"9a450002",
		16#0a77# => X"dc0f8800",
		16#0a78# => X"e2539002",
		16#0a79# => X"99e50000",
		16#0a7a# => X"a62fffff",
		16#0a7b# => X"e1ef2003",
		16#0a7c# => X"ba310048",
		16#0a7d# => X"bd520000",
		16#0a7e# => X"e1f17804",
		16#0a7f# => X"0fffffbe",
		16#0a80# => X"dc057800",
		16#0a81# => X"a8a20000",
		16#0a82# => X"84420000",
		16#0a83# => X"9d08ffff",
		16#0a84# => X"03ffffbc",
		16#0a85# => X"e1a01002",
		16#0a86# => X"0fffffc7",
		16#0a87# => X"bc220000",
		16#0a88# => X"03fffffa",
		16#0a89# => X"a8a20000",
		16#0a8a# => X"84620004",
		16#0a8b# => X"84c1000c",
		16#0a8c# => X"8c830001",
		16#0a8d# => X"e4243000",
		16#0a8e# => X"10000009",
		16#0a8f# => X"a9c20000",
		16#0a90# => X"03ffff85",
		16#0a91# => X"98630000",
		16#0a92# => X"848e0004",
		16#0a93# => X"8c840001",
		16#0a94# => X"e4242800",
		16#0a95# => X"0fffff7f",
		16#0a96# => X"15000000",
		16#0a97# => X"85ce0000",
		16#0a98# => X"bc0e0000",
		16#0a99# => X"0ffffff9",
		16#0a9a# => X"84a1000c",
		16#0a9b# => X"03ffff37",
		16#0a9c# => X"84820000",
		16#0a9d# => X"9d800000",
		16#0a9e# => X"ab8e0000",
		16#0a9f# => X"a90c0000",
		16#0aa0# => X"03fffed9",
		16#0aa1# => X"a96c0000",
		16#0aa2# => X"03ffff72",
		16#0aa3# => X"a9c20000",
		16#0aa4# => X"84500000",
		16#0aa5# => X"bc220000",
		16#0aa6# => X"0fffffb3",
		16#0aa7# => X"85610010",
		16#0aa8# => X"84700004",
		16#0aa9# => X"84810010",
		16#0aaa# => X"04001029",
		16#0aab# => X"98630000",
		16#0aac# => X"84420000",
		16#0aad# => X"bc220000",
		16#0aae# => X"13fffffa",
		16#0aaf# => X"d4015810",
		16#0ab0# => X"03ffffa9",
		16#0ab1# => X"85610010",
		16#0ab2# => X"b8a50010",
		16#0ab3# => X"d7e117f0",
		16#0ab4# => X"d7e187f8",
		16#0ab5# => X"a8440000",
		16#0ab6# => X"d7e14ffc",
		16#0ab7# => X"d7e177f4",
		16#0ab8# => X"9c800014",
		16#0ab9# => X"9c21fff0",
		16#0aba# => X"04001b12",
		16#0abb# => X"ba050090",
		16#0abc# => X"9c6bfffe",
		16#0abd# => X"9c800000",
		16#0abe# => X"b8e30003",
		16#0abf# => X"9ca00000",
		16#0ac0# => X"9d608080",
		16#0ac1# => X"e0e23800",
		16#0ac2# => X"d4022000",
		16#0ac3# => X"d4023804",
		16#0ac4# => X"b9e30002",
		16#0ac5# => X"9d020010",
		16#0ac6# => X"dc072802",
		16#0ac7# => X"dc075800",
		16#0ac8# => X"9c820008",
		16#0ac9# => X"e1e77800",
		16#0aca# => X"e4a74000",
		16#0acb# => X"10000006",
		16#0acc# => X"9ca70004",
		16#0acd# => X"9cc70008",
		16#0ace# => X"e4af3000",
		16#0acf# => X"0c0000a5",
		16#0ad0# => X"9dc00000",
		16#0ad1# => X"bc030000",
		16#0ad2# => X"10000023",
		16#0ad3# => X"a630ffff",
		16#0ad4# => X"85020000",
		16#0ad5# => X"00000018",
		16#0ad6# => X"9cc00000",
		16#0ad7# => X"a5a6ffff",
		16#0ad8# => X"e44f6000",
		16#0ad9# => X"e1cd8805",
		16#0ada# => X"a5ad0007",
		16#0adb# => X"0c000016",
		16#0adc# => X"a5ce000f",
		16#0add# => X"b9ce0003",
		16#0ade# => X"d4044000",
		16#0adf# => X"9d007fff",
		16#0ae0# => X"e1ae6804",
		16#0ae1# => X"d4042804",
		16#0ae2# => X"b9cd0008",
		16#0ae3# => X"d4022000",
		16#0ae4# => X"dc054002",
		16#0ae5# => X"e1ae6804",
		16#0ae6# => X"9cc60001",
		16#0ae7# => X"dc056800",
		16#0ae8# => X"a9040000",
		16#0ae9# => X"a8ac0000",
		16#0aea# => X"e4433000",
		16#0aeb# => X"0c00000a",
		16#0aec# => X"a88b0000",
		16#0aed# => X"9d640008",
		16#0aee# => X"e4475800",
		16#0aef# => X"13ffffe8",
		16#0af0# => X"9d850004",
		16#0af1# => X"9cc60001",
		16#0af2# => X"e4433000",
		16#0af3# => X"13fffffa",
		16#0af4# => X"85020000",
		16#0af5# => X"9c800005",
		16#0af6# => X"04001ad6",
		16#0af7# => X"85c20000",
		16#0af8# => X"9c800001",
		16#0af9# => X"00000008",
		16#0afa# => X"9c600002",
		16#0afb# => X"84ce0004",
		16#0afc# => X"dc062002",
		16#0afd# => X"9c840001",
		16#0afe# => X"9c630001",
		16#0aff# => X"a484ffff",
		16#0b00# => X"a9c50000",
		16#0b01# => X"a4e30007",
		16#0b02# => X"e0c48005",
		16#0b03# => X"b8e70008",
		16#0b04# => X"84ae0000",
		16#0b05# => X"9d03ffff",
		16#0b06# => X"e0c73004",
		16#0b07# => X"bc250000",
		16#0b08# => X"0c000008",
		16#0b09# => X"a4c63fff",
		16#0b0a# => X"e4685800",
		16#0b0b# => X"0ffffff0",
		16#0b0c# => X"15000000",
		16#0b0d# => X"84ee0004",
		16#0b0e# => X"03ffffef",
		16#0b0f# => X"dc073002",
		16#0b10# => X"bc020000",
		16#0b11# => X"10000034",
		16#0b12# => X"9cc00001",
		16#0b13# => X"9d600000",
		16#0b14# => X"a8a20000",
		16#0b15# => X"a8eb0000",
		16#0b16# => X"a9eb0000",
		16#0b17# => X"9def0001",
		16#0b18# => X"a8850000",
		16#0b19# => X"9c600000",
		16#0b1a# => X"84840000",
		16#0b1b# => X"bc240000",
		16#0b1c# => X"0c000005",
		16#0b1d# => X"9c630001",
		16#0b1e# => X"e5833000",
		16#0b1f# => X"13fffffb",
		16#0b20# => X"15000000",
		16#0b21# => X"a9850000",
		16#0b22# => X"a9060000",
		16#0b23# => X"a8a40000",
		16#0b24# => X"bd430000",
		16#0b25# => X"0c000011",
		16#0b26# => X"e1a02002",
		16#0b27# => X"e0856804",
		16#0b28# => X"bd640000",
		16#0b29# => X"0c000027",
		16#0b2a# => X"e0404002",
		16#0b2b# => X"a88c0000",
		16#0b2c# => X"9c63ffff",
		16#0b2d# => X"858c0000",
		16#0b2e# => X"bc070000",
		16#0b2f# => X"1000001e",
		16#0b30# => X"15000000",
		16#0b31# => X"d4072000",
		16#0b32# => X"a8e40000",
		16#0b33# => X"bd430000",
		16#0b34# => X"13fffff4",
		16#0b35# => X"e0856804",
		16#0b36# => X"e0856804",
		16#0b37# => X"bd640000",
		16#0b38# => X"0c000035",
		16#0b39# => X"bd480000",
		16#0b3a# => X"bc250000",
		16#0b3b# => X"13ffffdd",
		16#0b3c# => X"9def0001",
		16#0b3d# => X"9defffff",
		16#0b3e# => X"bc2f0001",
		16#0b3f# => X"0c000008",
		16#0b40# => X"d4072800",
		16#0b41# => X"a84b0000",
		16#0b42# => X"bc020000",
		16#0b43# => X"0fffffd0",
		16#0b44# => X"e0c63000",
		16#0b45# => X"d4021000",
		16#0b46# => X"a9620000",
		16#0b47# => X"9c210010",
		16#0b48# => X"8521fffc",
		16#0b49# => X"8441fff0",
		16#0b4a# => X"85c1fff4",
		16#0b4b# => X"44004800",
		16#0b4c# => X"8601fff8",
		16#0b4d# => X"a9640000",
		16#0b4e# => X"03ffffe5",
		16#0b4f# => X"a8e40000",
		16#0b50# => X"e0424004",
		16#0b51# => X"bd820000",
		16#0b52# => X"0fffffda",
		16#0b53# => X"a88c0000",
		16#0b54# => X"862c0004",
		16#0b55# => X"9dc0ff00",
		16#0b56# => X"9a710000",
		16#0b57# => X"a453ffff",
		16#0b58# => X"e2737003",
		16#0b59# => X"b8420048",
		16#0b5a# => X"84850004",
		16#0b5b# => X"9ab10002",
		16#0b5c# => X"e2629804",
		16#0b5d# => X"98440002",
		16#0b5e# => X"dc119800",
		16#0b5f# => X"e2751002",
		16#0b60# => X"9a240000",
		16#0b61# => X"a451ffff",
		16#0b62# => X"e2317003",
		16#0b63# => X"b8420048",
		16#0b64# => X"bd530000",
		16#0b65# => X"e2228804",
		16#0b66# => X"0fffffc5",
		16#0b67# => X"dc048800",
		16#0b68# => X"a8850000",
		16#0b69# => X"84a50000",
		16#0b6a# => X"9d08ffff",
		16#0b6b# => X"03ffffc3",
		16#0b6c# => X"e1a02802",
		16#0b6d# => X"0fffffce",
		16#0b6e# => X"bc250000",
		16#0b6f# => X"bc230000",
		16#0b70# => X"0ffffff8",
		16#0b71# => X"15000000",
		16#0b72# => X"03ffffb6",
		16#0b73# => X"e0856804",
		16#0b74# => X"d4042804",
		16#0b75# => X"d4047000",
		16#0b76# => X"d4022000",
		16#0b77# => X"9d607fff",
		16#0b78# => X"9c80ffff",
		16#0b79# => X"dc055802",
		16#0b7a# => X"dc052000",
		16#0b7b# => X"a8880000",
		16#0b7c# => X"03ffff55",
		16#0b7d# => X"a8a60000",
		16#0b7e# => X"85650000",
		16#0b7f# => X"d7e117fc",
		16#0b80# => X"9d8b0008",
		16#0b81# => X"e46c3800",
		16#0b82# => X"0c000006",
		16#0b83# => X"9c21fffc",
		16#0b84# => X"9d600000",
		16#0b85# => X"9c210004",
		16#0b86# => X"44004800",
		16#0b87# => X"8441fffc",
		16#0b88# => X"84e60000",
		16#0b89# => X"9da70004",
		16#0b8a# => X"e4a86800",
		16#0b8b# => X"13fffff9",
		16#0b8c# => X"15000000",
		16#0b8d# => X"d4056000",
		16#0b8e# => X"d40b3804",
		16#0b8f# => X"84e30000",
		16#0b90# => X"84a60000",
		16#0b91# => X"d40b3800",
		16#0b92# => X"9ca50004",
		16#0b93# => X"d4035800",
		16#0b94# => X"d4062800",
		16#0b95# => X"94440000",
		16#0b96# => X"94840002",
		16#0b97# => X"846b0004",
		16#0b98# => X"dc031000",
		16#0b99# => X"03ffffec",
		16#0b9a# => X"dc032002",
		16#0b9b# => X"85630000",
		16#0b9c# => X"d7e117fc",
		16#0b9d# => X"84cb0004",
		16#0b9e# => X"84ab0000",
		16#0b9f# => X"84830004",
		16#0ba0# => X"9c400000",
		16#0ba1# => X"9c21fffc",
		16#0ba2# => X"d4033004",
		16#0ba3# => X"d4032800",
		16#0ba4# => X"d40b1000",
		16#0ba5# => X"d40b2004",
		16#0ba6# => X"9c210004",
		16#0ba7# => X"44004800",
		16#0ba8# => X"8441fffc",
		16#0ba9# => X"84c40004",
		16#0baa# => X"84e40000",
		16#0bab# => X"84a30004",
		16#0bac# => X"d4033800",
		16#0bad# => X"d4033004",
		16#0bae# => X"d4042804",
		16#0baf# => X"d4041800",
		16#0bb0# => X"44004800",
		16#0bb1# => X"a9630000",
		16#0bb2# => X"98a40002",
		16#0bb3# => X"bd650000",
		16#0bb4# => X"0c000016",
		16#0bb5# => X"bc030000",
		16#0bb6# => X"10000012",
		16#0bb7# => X"a9630000",
		16#0bb8# => X"84830004",
		16#0bb9# => X"98840002",
		16#0bba# => X"e4042800",
		16#0bbb# => X"0c000009",
		16#0bbc# => X"15000000",
		16#0bbd# => X"0000000b",
		16#0bbe# => X"15000000",
		16#0bbf# => X"84830004",
		16#0bc0# => X"98840002",
		16#0bc1# => X"e4242800",
		16#0bc2# => X"0c000006",
		16#0bc3# => X"15000000",
		16#0bc4# => X"84630000",
		16#0bc5# => X"bc030000",
		16#0bc6# => X"0ffffff9",
		16#0bc7# => X"a9630000",
		16#0bc8# => X"44004800",
		16#0bc9# => X"15000000",
		16#0bca# => X"13fffffe",
		16#0bcb# => X"a9630000",
		16#0bcc# => X"84c30004",
		16#0bcd# => X"98a40000",
		16#0bce# => X"8c860001",
		16#0bcf# => X"e4242800",
		16#0bd0# => X"10000009",
		16#0bd1# => X"15000000",
		16#0bd2# => X"03fffff6",
		16#0bd3# => X"15000000",
		16#0bd4# => X"84830004",
		16#0bd5# => X"8c840001",
		16#0bd6# => X"e4242800",
		16#0bd7# => X"0ffffff1",
		16#0bd8# => X"a9630000",
		16#0bd9# => X"84630000",
		16#0bda# => X"bc030000",
		16#0bdb# => X"0ffffff9",
		16#0bdc# => X"15000000",
		16#0bdd# => X"44004800",
		16#0bde# => X"a9630000",
		16#0bdf# => X"bc030000",
		16#0be0# => X"0c000005",
		16#0be1# => X"9ca00000",
		16#0be2# => X"00000009",
		16#0be3# => X"a9630000",
		16#0be4# => X"a8640000",
		16#0be5# => X"84830000",
		16#0be6# => X"d4032800",
		16#0be7# => X"bc240000",
		16#0be8# => X"13fffffc",
		16#0be9# => X"a8a30000",
		16#0bea# => X"a9630000",
		16#0beb# => X"44004800",
		16#0bec# => X"15000000",
		16#0bed# => X"d7e187dc",
		16#0bee# => X"d7e1e7f4",
		16#0bef# => X"d7e1f7f8",
		16#0bf0# => X"d7e14ffc",
		16#0bf1# => X"d7e117d4",
		16#0bf2# => X"d7e177d8",
		16#0bf3# => X"d7e197e0",
		16#0bf4# => X"d7e1a7e4",
		16#0bf5# => X"d7e1b7e8",
		16#0bf6# => X"d7e1c7ec",
		16#0bf7# => X"d7e1d7f0",
		16#0bf8# => X"9c21ffd0",
		16#0bf9# => X"ab830000",
		16#0bfa# => X"d4012000",
		16#0bfb# => X"abc50000",
		16#0bfc# => X"bc1c0000",
		16#0bfd# => X"10000049",
		16#0bfe# => X"9e000001",
		16#0bff# => X"9f400000",
		16#0c00# => X"aa9c0000",
		16#0c01# => X"aa5a0000",
		16#0c02# => X"ab9a0000",
		16#0c03# => X"9f5a0001",
		16#0c04# => X"a8540000",
		16#0c05# => X"9dc00000",
		16#0c06# => X"84420000",
		16#0c07# => X"bc220000",
		16#0c08# => X"0c000005",
		16#0c09# => X"9dce0001",
		16#0c0a# => X"e5507000",
		16#0c0b# => X"13fffffb",
		16#0c0c# => X"15000000",
		16#0c0d# => X"aad00000",
		16#0c0e# => X"bc2e0000",
		16#0c0f# => X"0c000011",
		16#0c10# => X"e3001002",
		16#0c11# => X"e0c2c004",
		16#0c12# => X"bd660000",
		16#0c13# => X"0c000018",
		16#0c14# => X"e060b002",
		16#0c15# => X"a8d40000",
		16#0c16# => X"9dceffff",
		16#0c17# => X"86940000",
		16#0c18# => X"bc120000",
		16#0c19# => X"1000000f",
		16#0c1a# => X"15000000",
		16#0c1b# => X"d4123000",
		16#0c1c# => X"aa460000",
		16#0c1d# => X"bc2e0000",
		16#0c1e# => X"13fffff4",
		16#0c1f# => X"e0c2c004",
		16#0c20# => X"e302c004",
		16#0c21# => X"bd780000",
		16#0c22# => X"0c00001a",
		16#0c23# => X"bc220000",
		16#0c24# => X"0c00001d",
		16#0c25# => X"bc3a0001",
		16#0c26# => X"03ffffdd",
		16#0c27# => X"aa820000",
		16#0c28# => X"ab860000",
		16#0c29# => X"03fffff4",
		16#0c2a# => X"aa460000",
		16#0c2b# => X"e063b004",
		16#0c2c# => X"bd830000",
		16#0c2d# => X"0fffffe9",
		16#0c2e# => X"a8d40000",
		16#0c2f# => X"84740004",
		16#0c30# => X"84820004",
		16#0c31# => X"84c10000",
		16#0c32# => X"48003000",
		16#0c33# => X"a8be0000",
		16#0c34# => X"bd4b0000",
		16#0c35# => X"0fffffe0",
		16#0c36# => X"15000000",
		16#0c37# => X"a8c20000",
		16#0c38# => X"84420000",
		16#0c39# => X"9ed6ffff",
		16#0c3a# => X"03ffffde",
		16#0c3b# => X"e3001002",
		16#0c3c# => X"bd560000",
		16#0c3d# => X"13fffffa",
		16#0c3e# => X"bc220000",
		16#0c3f# => X"13ffffe7",
		16#0c40# => X"bc3a0001",
		16#0c41# => X"0c000006",
		16#0c42# => X"d4121000",
		16#0c43# => X"bc1c0000",
		16#0c44# => X"0fffffbb",
		16#0c45# => X"e2108000",
		16#0c46# => X"d41ce000",
		16#0c47# => X"9c210030",
		16#0c48# => X"a97c0000",
		16#0c49# => X"8521fffc",
		16#0c4a# => X"8441ffd4",
		16#0c4b# => X"85c1ffd8",
		16#0c4c# => X"8601ffdc",
		16#0c4d# => X"8641ffe0",
		16#0c4e# => X"8681ffe4",
		16#0c4f# => X"86c1ffe8",
		16#0c50# => X"8701ffec",
		16#0c51# => X"8741fff0",
		16#0c52# => X"8781fff4",
		16#0c53# => X"44004800",
		16#0c54# => X"87c1fff8",
		16#0c55# => X"d7e117f0",
		16#0c56# => X"d7e187f8",
		16#0c57# => X"a8430000",
		16#0c58# => X"8603001c",
		16#0c59# => X"9c600000",
		16#0c5a# => X"d7e14ffc",
		16#0c5b# => X"d7e177f4",
		16#0c5c# => X"dc021838",
		16#0c5d# => X"dc02183a",
		16#0c5e# => X"dc02183c",
		16#0c5f# => X"dc02183e",
		16#0c60# => X"bc100000",
		16#0c61# => X"10000018",
		16#0c62# => X"9c21fff0",
		16#0c63# => X"9dc00000",
		16#0c64# => X"9c800001",
		16#0c65# => X"07fffcba",
		16#0c66# => X"a8620000",
		16#0c67# => X"94820038",
		16#0c68# => X"04000c53",
		16#0c69# => X"a86b0000",
		16#0c6a# => X"9c80ffff",
		16#0c6b# => X"a8620000",
		16#0c6c# => X"07fffcb3",
		16#0c6d# => X"dc025838",
		16#0c6e# => X"94820038",
		16#0c6f# => X"04000c4c",
		16#0c70# => X"a86b0000",
		16#0c71# => X"dc025838",
		16#0c72# => X"bc2e0000",
		16#0c73# => X"10000003",
		16#0c74# => X"9dce0001",
		16#0c75# => X"dc02583a",
		16#0c76# => X"e4507000",
		16#0c77# => X"13ffffee",
		16#0c78# => X"9c800001",
		16#0c79# => X"9c210010",
		16#0c7a# => X"9d600000",
		16#0c7b# => X"8521fffc",
		16#0c7c# => X"8441fff0",
		16#0c7d# => X"85c1fff4",
		16#0c7e# => X"44004800",
		16#0c7f# => X"8601fff8",
		16#0c80# => X"d7e14ffc",
		16#0c81# => X"d7e117d4",
		16#0c82# => X"d7e177d8",
		16#0c83# => X"d7e187dc",
		16#0c84# => X"d7e197e0",
		16#0c85# => X"d7e1a7e4",
		16#0c86# => X"d7e1b7e8",
		16#0c87# => X"d7e1c7ec",
		16#0c88# => X"d7e1d7f0",
		16#0c89# => X"d7e1e7f4",
		16#0c8a# => X"d7e1f7f8",
		16#0c8b# => X"9c21fd54",
		16#0c8c# => X"a8a40000",
		16#0c8d# => X"d401181c",
		16#0c8e# => X"9c81001c",
		16#0c8f# => X"04000f5e",
		16#0c90# => X"9c610064",
		16#0c91# => X"04000ba2",
		16#0c92# => X"9c600001",
		16#0c93# => X"9c600002",
		16#0c94# => X"04000b9f",
		16#0c95# => X"dc015820",
		16#0c96# => X"9c600003",
		16#0c97# => X"04000b9c",
		16#0c98# => X"dc015822",
		16#0c99# => X"9c600004",
		16#0c9a# => X"04000b99",
		16#0c9b# => X"dc015824",
		16#0c9c# => X"9c600005",
		16#0c9d# => X"04000b96",
		16#0c9e# => X"d401583c",
		16#0c9f# => X"bc2b0000",
		16#0ca0# => X"10000004",
		16#0ca1# => X"d4015840",
		16#0ca2# => X"9c400007",
		16#0ca3# => X"d4011040",
		16#0ca4# => X"84410020",
		16#0ca5# => X"bc220000",
		16#0ca6# => X"10000305",
		16#0ca7# => X"18600001",
		16#0ca8# => X"98610024",
		16#0ca9# => X"bc230000",
		16#0caa# => X"0c0002fc",
		16#0cab# => X"18600001",
		16#0cac# => X"04000b87",
		16#0cad# => X"9c600007",
		16#0cae# => X"b84b0010",
		16#0caf# => X"b8420090",
		16#0cb0# => X"bc220000",
		16#0cb1# => X"1000030b",
		16#0cb2# => X"15000000",
		16#0cb3# => X"9c4007d0",
		16#0cb4# => X"d4011038",
		16#0cb5# => X"a8620000",
		16#0cb6# => X"04000ed3",
		16#0cb7# => X"9c400000",
		16#0cb8# => X"9c600007",
		16#0cb9# => X"dc011060",
		16#0cba# => X"04000b79",
		16#0cbb# => X"d4015828",
		16#0cbc# => X"b84b0010",
		16#0cbd# => X"b8420090",
		16#0cbe# => X"bc220000",
		16#0cbf# => X"10000305",
		16#0cc0# => X"15000000",
		16#0cc1# => X"9c4007d0",
		16#0cc2# => X"d4011084",
		16#0cc3# => X"04000ec6",
		16#0cc4# => X"a8620000",
		16#0cc5# => X"94410020",
		16#0cc6# => X"dc01106c",
		16#0cc7# => X"94410022",
		16#0cc8# => X"dc01106e",
		16#0cc9# => X"94410024",
		16#0cca# => X"dc011070",
		16#0ccb# => X"9c400000",
		16#0ccc# => X"9c600007",
		16#0ccd# => X"dc0110ac",
		16#0cce# => X"84410040",
		16#0ccf# => X"d4015874",
		16#0cd0# => X"04000b63",
		16#0cd1# => X"d401108c",
		16#0cd2# => X"b84b0010",
		16#0cd3# => X"b8420090",
		16#0cd4# => X"bc220000",
		16#0cd5# => X"100002ed",
		16#0cd6# => X"15000000",
		16#0cd7# => X"9c4007d0",
		16#0cd8# => X"d40110d0",
		16#0cd9# => X"04000eb0",
		16#0cda# => X"a8620000",
		16#0cdb# => X"94410020",
		16#0cdc# => X"dc0110b8",
		16#0cdd# => X"94410022",
		16#0cde# => X"dc0110ba",
		16#0cdf# => X"94410024",
		16#0ce0# => X"dc0110bc",
		16#0ce1# => X"9c400000",
		16#0ce2# => X"9c600007",
		16#0ce3# => X"dc0110f8",
		16#0ce4# => X"84410040",
		16#0ce5# => X"d40158c0",
		16#0ce6# => X"04000b4d",
		16#0ce7# => X"d40110d8",
		16#0ce8# => X"b84b0010",
		16#0ce9# => X"b8420090",
		16#0cea# => X"bc220000",
		16#0ceb# => X"100002e1",
		16#0cec# => X"15000000",
		16#0ced# => X"9c4007d0",
		16#0cee# => X"d401111c",
		16#0cef# => X"04000e9a",
		16#0cf0# => X"a8620000",
		16#0cf1# => X"94410020",
		16#0cf2# => X"dc011104",
		16#0cf3# => X"94410022",
		16#0cf4# => X"dc011106",
		16#0cf5# => X"94410024",
		16#0cf6# => X"dc011108",
		16#0cf7# => X"9c400000",
		16#0cf8# => X"9c600007",
		16#0cf9# => X"dc011144",
		16#0cfa# => X"84410040",
		16#0cfb# => X"d401590c",
		16#0cfc# => X"04000b37",
		16#0cfd# => X"d4011124",
		16#0cfe# => X"b84b0010",
		16#0cff# => X"b8420090",
		16#0d00# => X"bc220000",
		16#0d01# => X"100002c9",
		16#0d02# => X"15000000",
		16#0d03# => X"9c4007d0",
		16#0d04# => X"d4011168",
		16#0d05# => X"04000e84",
		16#0d06# => X"a8620000",
		16#0d07# => X"94410020",
		16#0d08# => X"dc011150",
		16#0d09# => X"94410022",
		16#0d0a# => X"dc011152",
		16#0d0b# => X"94410024",
		16#0d0c# => X"dc011154",
		16#0d0d# => X"9c400000",
		16#0d0e# => X"9c600007",
		16#0d0f# => X"dc011190",
		16#0d10# => X"84410040",
		16#0d11# => X"d4015958",
		16#0d12# => X"04000b21",
		16#0d13# => X"d4011170",
		16#0d14# => X"b84b0010",
		16#0d15# => X"b8420090",
		16#0d16# => X"bc220000",
		16#0d17# => X"100002b1",
		16#0d18# => X"15000000",
		16#0d19# => X"9c4007d0",
		16#0d1a# => X"d40111b4",
		16#0d1b# => X"04000e6e",
		16#0d1c# => X"a8620000",
		16#0d1d# => X"94410020",
		16#0d1e# => X"dc01119c",
		16#0d1f# => X"94410022",
		16#0d20# => X"dc01119e",
		16#0d21# => X"94410024",
		16#0d22# => X"dc0111a0",
		16#0d23# => X"9c400000",
		16#0d24# => X"9c600007",
		16#0d25# => X"dc0111dc",
		16#0d26# => X"84410040",
		16#0d27# => X"d40159a4",
		16#0d28# => X"04000b0b",
		16#0d29# => X"d40111bc",
		16#0d2a# => X"b84b0010",
		16#0d2b# => X"b8420090",
		16#0d2c# => X"bc220000",
		16#0d2d# => X"10000299",
		16#0d2e# => X"15000000",
		16#0d2f# => X"9c4007d0",
		16#0d30# => X"d4011200",
		16#0d31# => X"04000e58",
		16#0d32# => X"a8620000",
		16#0d33# => X"94410020",
		16#0d34# => X"dc0111e8",
		16#0d35# => X"94410022",
		16#0d36# => X"dc0111ea",
		16#0d37# => X"94410024",
		16#0d38# => X"dc0111ec",
		16#0d39# => X"9c400000",
		16#0d3a# => X"9c600007",
		16#0d3b# => X"dc011228",
		16#0d3c# => X"84410040",
		16#0d3d# => X"d40159f0",
		16#0d3e# => X"04000af5",
		16#0d3f# => X"d4011208",
		16#0d40# => X"b84b0010",
		16#0d41# => X"b8420090",
		16#0d42# => X"bc020000",
		16#0d43# => X"0c000004",
		16#0d44# => X"a8620000",
		16#0d45# => X"9c4007d0",
		16#0d46# => X"a8620000",
		16#0d47# => X"04000e42",
		16#0d48# => X"d401124c",
		16#0d49# => X"94610020",
		16#0d4a# => X"dc011a34",
		16#0d4b# => X"94610022",
		16#0d4c# => X"dc011a36",
		16#0d4d# => X"94610024",
		16#0d4e# => X"84410040",
		16#0d4f# => X"dc011a38",
		16#0d50# => X"9c600000",
		16#0d51# => X"a5c20001",
		16#0d52# => X"d4015a3c",
		16#0d53# => X"dc011a74",
		16#0d54# => X"bc0e0000",
		16#0d55# => X"10000003",
		16#0d56# => X"d4011254",
		16#0d57# => X"9dc00001",
		16#0d58# => X"9c8e0001",
		16#0d59# => X"a4620002",
		16#0d5a# => X"bc030000",
		16#0d5b# => X"10000003",
		16#0d5c# => X"a484ffff",
		16#0d5d# => X"a9c40000",
		16#0d5e# => X"9c8e0001",
		16#0d5f# => X"a4620004",
		16#0d60# => X"bc030000",
		16#0d61# => X"10000003",
		16#0d62# => X"a484ffff",
		16#0d63# => X"a9c40000",
		16#0d64# => X"a5ceffff",
		16#0d65# => X"84610038",
		16#0d66# => X"04001866",
		16#0d67# => X"a88e0000",
		16#0d68# => X"84610084",
		16#0d69# => X"a88e0000",
		16#0d6a# => X"aa0b0000",
		16#0d6b# => X"04001861",
		16#0d6c# => X"d4015838",
		16#0d6d# => X"846100d0",
		16#0d6e# => X"a88e0000",
		16#0d6f# => X"0400185d",
		16#0d70# => X"d4015884",
		16#0d71# => X"8461011c",
		16#0d72# => X"a88e0000",
		16#0d73# => X"04001859",
		16#0d74# => X"d40158d0",
		16#0d75# => X"84610168",
		16#0d76# => X"a88e0000",
		16#0d77# => X"04001855",
		16#0d78# => X"d401591c",
		16#0d79# => X"846101b4",
		16#0d7a# => X"a88e0000",
		16#0d7b# => X"04001851",
		16#0d7c# => X"d4015968",
		16#0d7d# => X"84610200",
		16#0d7e# => X"a88e0000",
		16#0d7f# => X"0400184d",
		16#0d80# => X"d40159b4",
		16#0d81# => X"8461024c",
		16#0d82# => X"a88e0000",
		16#0d83# => X"04001849",
		16#0d84# => X"d4015a00",
		16#0d85# => X"a4820001",
		16#0d86# => X"bc040000",
		16#0d87# => X"10000013",
		16#0d88# => X"d4015a4c",
		16#0d89# => X"84610028",
		16#0d8a# => X"9c800001",
		16#0d8b# => X"d401182c",
		16#0d8c# => X"84610074",
		16#0d8d# => X"d4011878",
		16#0d8e# => X"846100c0",
		16#0d8f# => X"d40118c4",
		16#0d90# => X"8461010c",
		16#0d91# => X"d4011910",
		16#0d92# => X"84610158",
		16#0d93# => X"d401195c",
		16#0d94# => X"846101a4",
		16#0d95# => X"d40119a8",
		16#0d96# => X"846101f0",
		16#0d97# => X"d40119f4",
		16#0d98# => X"8461023c",
		16#0d99# => X"d4011a40",
		16#0d9a# => X"a4620002",
		16#0d9b# => X"bc030000",
		16#0d9c# => X"1000001e",
		16#0d9d# => X"a4620004",
		16#0d9e# => X"e0a48306",
		16#0d9f# => X"85a10028",
		16#0da0# => X"85810074",
		16#0da1# => X"856100c0",
		16#0da2# => X"8501010c",
		16#0da3# => X"84e10158",
		16#0da4# => X"84c101a4",
		16#0da5# => X"846101f0",
		16#0da6# => X"85c1023c",
		16#0da7# => X"e1ad2800",
		16#0da8# => X"e18c2800",
		16#0da9# => X"e16b2800",
		16#0daa# => X"e1082800",
		16#0dab# => X"e0e72800",
		16#0dac# => X"e0c62800",
		16#0dad# => X"e0632800",
		16#0dae# => X"9c840001",
		16#0daf# => X"e0ae2800",
		16#0db0# => X"d4016830",
		16#0db1# => X"d401607c",
		16#0db2# => X"d40158c8",
		16#0db3# => X"d4014114",
		16#0db4# => X"d4013960",
		16#0db5# => X"d40131ac",
		16#0db6# => X"d40119f8",
		16#0db7# => X"d4012a44",
		16#0db8# => X"a484ffff",
		16#0db9# => X"a4620004",
		16#0dba# => X"bc030000",
		16#0dbb# => X"1000001c",
		16#0dbc# => X"a4620001",
		16#0dbd# => X"e0848306",
		16#0dbe# => X"85810028",
		16#0dbf# => X"85610074",
		16#0dc0# => X"850100c0",
		16#0dc1# => X"84e1010c",
		16#0dc2# => X"84c10158",
		16#0dc3# => X"84a101a4",
		16#0dc4# => X"846101f0",
		16#0dc5# => X"85a1023c",
		16#0dc6# => X"e18c2000",
		16#0dc7# => X"e16b2000",
		16#0dc8# => X"e1082000",
		16#0dc9# => X"e0e72000",
		16#0dca# => X"e0c62000",
		16#0dcb# => X"e0a52000",
		16#0dcc# => X"e0632000",
		16#0dcd# => X"e08d2000",
		16#0dce# => X"d4016034",
		16#0dcf# => X"d4015880",
		16#0dd0# => X"d40140cc",
		16#0dd1# => X"d4013918",
		16#0dd2# => X"d4013164",
		16#0dd3# => X"d40129b0",
		16#0dd4# => X"d40119fc",
		16#0dd5# => X"d4012248",
		16#0dd6# => X"a4620001",
		16#0dd7# => X"bc030000",
		16#0dd8# => X"0c0002d9",
		16#0dd9# => X"84610038",
		16#0dda# => X"a4620002",
		16#0ddb# => X"bc030000",
		16#0ddc# => X"0c00024f",
		16#0ddd# => X"a4420004",
		16#0dde# => X"bc020000",
		16#0ddf# => X"0c000259",
		16#0de0# => X"8441008c",
		16#0de1# => X"a4620001",
		16#0de2# => X"bc030000",
		16#0de3# => X"0c00025e",
		16#0de4# => X"a4620002",
		16#0de5# => X"bc030000",
		16#0de6# => X"0c000264",
		16#0de7# => X"15000000",
		16#0de8# => X"a4420004",
		16#0de9# => X"bc020000",
		16#0dea# => X"0c00026d",
		16#0deb# => X"844100d8",
		16#0dec# => X"a4620001",
		16#0ded# => X"bc030000",
		16#0dee# => X"0c000272",
		16#0def# => X"a4620002",
		16#0df0# => X"bc030000",
		16#0df1# => X"0c000278",
		16#0df2# => X"15000000",
		16#0df3# => X"a4420004",
		16#0df4# => X"bc020000",
		16#0df5# => X"0c000281",
		16#0df6# => X"84410124",
		16#0df7# => X"a4620001",
		16#0df8# => X"bc030000",
		16#0df9# => X"0c000286",
		16#0dfa# => X"a4620002",
		16#0dfb# => X"bc030000",
		16#0dfc# => X"0c00028c",
		16#0dfd# => X"15000000",
		16#0dfe# => X"a4420004",
		16#0dff# => X"bc020000",
		16#0e00# => X"0c000295",
		16#0e01# => X"84410170",
		16#0e02# => X"a4620001",
		16#0e03# => X"bc030000",
		16#0e04# => X"0c00029a",
		16#0e05# => X"a4620002",
		16#0e06# => X"bc030000",
		16#0e07# => X"0c0002a0",
		16#0e08# => X"15000000",
		16#0e09# => X"a4420004",
		16#0e0a# => X"bc020000",
		16#0e0b# => X"0c00021b",
		16#0e0c# => X"84610038",
		16#0e0d# => X"844101bc",
		16#0e0e# => X"a4620001",
		16#0e0f# => X"bc030000",
		16#0e10# => X"0c000210",
		16#0e11# => X"84610038",
		16#0e12# => X"a4620002",
		16#0e13# => X"bc030000",
		16#0e14# => X"0c000203",
		16#0e15# => X"84610038",
		16#0e16# => X"a4420004",
		16#0e17# => X"bc020000",
		16#0e18# => X"0c0001fa",
		16#0e19# => X"84610038",
		16#0e1a# => X"84410208",
		16#0e1b# => X"a4620001",
		16#0e1c# => X"bc030000",
		16#0e1d# => X"0c0001ef",
		16#0e1e# => X"84610038",
		16#0e1f# => X"a4620002",
		16#0e20# => X"bc030000",
		16#0e21# => X"0c0001e2",
		16#0e22# => X"84610038",
		16#0e23# => X"a4420004",
		16#0e24# => X"bc020000",
		16#0e25# => X"0c0001d9",
		16#0e26# => X"84610038",
		16#0e27# => X"84410254",
		16#0e28# => X"a4620001",
		16#0e29# => X"bc030000",
		16#0e2a# => X"0c0001b9",
		16#0e2b# => X"a4620002",
		16#0e2c# => X"bc030000",
		16#0e2d# => X"0c0001bf",
		16#0e2e# => X"15000000",
		16#0e2f# => X"a4420004",
		16#0e30# => X"bc020000",
		16#0e31# => X"0c0001c8",
		16#0e32# => X"98810234",
		16#0e33# => X"8441003c",
		16#0e34# => X"bc220000",
		16#0e35# => X"10000046",
		16#0e36# => X"1a400001",
		16#0e37# => X"9c400001",
		16#0e38# => X"aa528360",
		16#0e39# => X"9dc10020",
		16#0e3a# => X"b8820003",
		16#0e3b# => X"e0421000",
		16#0e3c# => X"e0422000",
		16#0e3d# => X"d401103c",
		16#0e3e# => X"04000d71",
		16#0e3f# => X"9c400000",
		16#0e40# => X"8601003c",
		16#0e41# => X"dc011058",
		16#0e42# => X"dc01105a",
		16#0e43# => X"dc01105c",
		16#0e44# => X"bc100000",
		16#0e45# => X"10000018",
		16#0e46# => X"dc01105e",
		16#0e47# => X"9c400000",
		16#0e48# => X"9c800001",
		16#0e49# => X"07fffad6",
		16#0e4a# => X"a86e0000",
		16#0e4b# => X"94810058",
		16#0e4c# => X"04000a6f",
		16#0e4d# => X"a86b0000",
		16#0e4e# => X"9c80ffff",
		16#0e4f# => X"a86e0000",
		16#0e50# => X"07fffacf",
		16#0e51# => X"dc015858",
		16#0e52# => X"94810058",
		16#0e53# => X"04000a68",
		16#0e54# => X"a86b0000",
		16#0e55# => X"dc015858",
		16#0e56# => X"bc220000",
		16#0e57# => X"10000003",
		16#0e58# => X"9c420001",
		16#0e59# => X"dc01585a",
		16#0e5a# => X"e4501000",
		16#0e5b# => X"13ffffee",
		16#0e5c# => X"9c800001",
		16#0e5d# => X"04000d6a",
		16#0e5e# => X"15000000",
		16#0e5f# => X"04000d72",
		16#0e60# => X"15000000",
		16#0e61# => X"04000d78",
		16#0e62# => X"a86b0000",
		16#0e63# => X"84b20000",
		16#0e64# => X"84d20004",
		16#0e65# => X"d4015810",
		16#0e66# => X"d4016014",
		16#0e67# => X"e06b0004",
		16#0e68# => X"e08c0004",
		16#0e69# => X"0400212e",
		16#0e6a# => X"15000000",
		16#0e6b# => X"bd8b0000",
		16#0e6c# => X"13ffffce",
		16#0e6d# => X"8441003c",
		16#0e6e# => X"84610010",
		16#0e6f# => X"84810014",
		16#0e70# => X"040017b4",
		16#0e71# => X"9c40000b",
		16#0e72# => X"bc0b0000",
		16#0e73# => X"10000005",
		16#0e74# => X"9c60000a",
		16#0e75# => X"04001757",
		16#0e76# => X"a88b0000",
		16#0e77# => X"9c4b0001",
		16#0e78# => X"8461003c",
		16#0e79# => X"e0431306",
		16#0e7a# => X"d401103c",
		16#0e7b# => X"04000d34",
		16#0e7c# => X"18400001",
		16#0e7d# => X"a842ade0",
		16#0e7e# => X"84620000",
		16#0e7f# => X"bca30008",
		16#0e80# => X"1000013e",
		16#0e81# => X"bc230000",
		16#0e82# => X"9c600008",
		16#0e83# => X"d4021800",
		16#0e84# => X"9c800000",
		16#0e85# => X"9e010020",
		16#0e86# => X"a9c40000",
		16#0e87# => X"9e40004c",
		16#0e88# => X"e0849306",
		16#0e89# => X"e0ae9306",
		16#0e8a# => X"9c610280",
		16#0e8b# => X"9dce0001",
		16#0e8c# => X"e0a32800",
		16#0e8d# => X"e0702000",
		16#0e8e# => X"8481003c",
		16#0e8f# => X"a5ceffff",
		16#0e90# => X"d7e525bc",
		16#0e91# => X"84810040",
		16#0e92# => X"04000db8",
		16#0e93# => X"d7e525c0",
		16#0e94# => X"84a20000",
		16#0e95# => X"e48e2800",
		16#0e96# => X"13fffff2",
		16#0e97# => X"a88e0000",
		16#0e98# => X"bc050000",
		16#0e99# => X"1000000e",
		16#0e9a# => X"15000000",
		16#0e9b# => X"9c800000",
		16#0e9c# => X"9e40004c",
		16#0e9d# => X"a9c40000",
		16#0e9e# => X"e0849306",
		16#0e9f# => X"e0702000",
		16#0ea0# => X"04000df3",
		16#0ea1# => X"9dce0001",
		16#0ea2# => X"a5ceffff",
		16#0ea3# => X"84a20000",
		16#0ea4# => X"e48e2800",
		16#0ea5# => X"13fffff9",
		16#0ea6# => X"a88e0000",
		16#0ea7# => X"04000d20",
		16#0ea8# => X"15000000",
		16#0ea9# => X"04000d28",
		16#0eaa# => X"15000000",
		16#0eab# => X"98610020",
		16#0eac# => X"9c800000",
		16#0ead# => X"04000c26",
		16#0eae# => X"ab4b0000",
		16#0eaf# => X"98610022",
		16#0eb0# => X"04000c23",
		16#0eb1# => X"a88b0000",
		16#0eb2# => X"98610024",
		16#0eb3# => X"04000c20",
		16#0eb4# => X"a88b0000",
		16#0eb5# => X"9861003a",
		16#0eb6# => X"04000c1d",
		16#0eb7# => X"a88b0000",
		16#0eb8# => X"bc0b7b05",
		16#0eb9# => X"10000454",
		16#0eba# => X"aacb0000",
		16#0ebb# => X"bc4b7b05",
		16#0ebc# => X"0c000112",
		16#0ebd# => X"bc0b18f2",
		16#0ebe# => X"a8608a02",
		16#0ebf# => X"e40b1800",
		16#0ec0# => X"1000045e",
		16#0ec1# => X"a860e9f5",
		16#0ec2# => X"e40b1800",
		16#0ec3# => X"100001f4",
		16#0ec4# => X"9c60ffff",
		16#0ec5# => X"aa40ffff",
		16#0ec6# => X"d4011818",
		16#0ec7# => X"04000cc0",
		16#0ec8# => X"15000000",
		16#0ec9# => X"040016d0",
		16#0eca# => X"e24b9000",
		16#0ecb# => X"ba520010",
		16#0ecc# => X"bc0b0000",
		16#0ecd# => X"0c00027f",
		16#0ece# => X"ba520090",
		16#0ecf# => X"040016ca",
		16#0ed0# => X"15000000",
		16#0ed1# => X"18600001",
		16#0ed2# => X"d4015800",
		16#0ed3# => X"040026ab",
		16#0ed4# => X"a8637ebc",
		16#0ed5# => X"18600001",
		16#0ed6# => X"84810038",
		16#0ed7# => X"a8638033",
		16#0ed8# => X"040026a6",
		16#0ed9# => X"d4012000",
		16#0eda# => X"040016bf",
		16#0edb# => X"15000000",
		16#0edc# => X"bc0b0000",
		16#0edd# => X"0c000401",
		16#0ede# => X"15000000",
		16#0edf# => X"040016ba",
		16#0ee0# => X"15000000",
		16#0ee1# => X"18600001",
		16#0ee2# => X"d4015800",
		16#0ee3# => X"0400269b",
		16#0ee4# => X"a8637ebc",
		16#0ee5# => X"18600001",
		16#0ee6# => X"d401d000",
		16#0ee7# => X"04002697",
		16#0ee8# => X"a863804b",
		16#0ee9# => X"040016b0",
		16#0eea# => X"15000000",
		16#0eeb# => X"bc0b0000",
		16#0eec# => X"0c0003ec",
		16#0eed# => X"15000000",
		16#0eee# => X"040016ab",
		16#0eef# => X"15000000",
		16#0ef0# => X"18600001",
		16#0ef1# => X"d4015800",
		16#0ef2# => X"0400268c",
		16#0ef3# => X"a8637ebc",
		16#0ef4# => X"04000ce5",
		16#0ef5# => X"a87a0000",
		16#0ef6# => X"18600001",
		16#0ef7# => X"d4015800",
		16#0ef8# => X"d4016004",
		16#0ef9# => X"04002685",
		16#0efa# => X"a8638063",
		16#0efb# => X"04000cde",
		16#0efc# => X"a87a0000",
		16#0efd# => X"18a00001",
		16#0efe# => X"e06b0004",
		16#0eff# => X"e08c0004",
		16#0f00# => X"a8a58368",
		16#0f01# => X"84c50004",
		16#0f02# => X"84a50000",
		16#0f03# => X"04002058",
		16#0f04# => X"15000000",
		16#0f05# => X"bd4b0000",
		16#0f06# => X"100003b2",
		16#0f07# => X"15000000",
		16#0f08# => X"04000cd1",
		16#0f09# => X"a87a0000",
		16#0f0a# => X"18a00001",
		16#0f0b# => X"e06b0004",
		16#0f0c# => X"e08c0004",
		16#0f0d# => X"a8a58370",
		16#0f0e# => X"84c50004",
		16#0f0f# => X"84a50000",
		16#0f10# => X"04002087",
		16#0f11# => X"15000000",
		16#0f12# => X"bd8b0000",
		16#0f13# => X"10000393",
		16#0f14# => X"15000000",
		16#0f15# => X"04001684",
		16#0f16# => X"15000000",
		16#0f17# => X"bc0b0000",
		16#0f18# => X"0c000388",
		16#0f19# => X"15000000",
		16#0f1a# => X"0400167f",
		16#0f1b# => X"15000000",
		16#0f1c# => X"18600001",
		16#0f1d# => X"d4015800",
		16#0f1e# => X"04002660",
		16#0f1f# => X"a8637ebc",
		16#0f20# => X"84a20000",
		16#0f21# => X"8481003c",
		16#0f22# => X"18600001",
		16#0f23# => X"e0852306",
		16#0f24# => X"a86380ce",
		16#0f25# => X"04002659",
		16#0f26# => X"d4012000",
		16#0f27# => X"04001672",
		16#0f28# => X"15000000",
		16#0f29# => X"bc0b0000",
		16#0f2a# => X"0c000370",
		16#0f2b# => X"15000000",
		16#0f2c# => X"0400166d",
		16#0f2d# => X"1bc00001",
		16#0f2e# => X"18600001",
		16#0f2f# => X"d4015800",
		16#0f30# => X"0400264e",
		16#0f31# => X"a8637ebc",
		16#0f32# => X"18600001",
		16#0f33# => X"abde80fd",
		16#0f34# => X"a86380e6",
		16#0f35# => X"04002649",
		16#0f36# => X"d401f000",
		16#0f37# => X"04001662",
		16#0f38# => X"15000000",
		16#0f39# => X"bc0b0000",
		16#0f3a# => X"0c00035a",
		16#0f3b# => X"15000000",
		16#0f3c# => X"0400165d",
		16#0f3d# => X"1b800001",
		16#0f3e# => X"18600001",
		16#0f3f# => X"d4015800",
		16#0f40# => X"0400263e",
		16#0f41# => X"a8637ebc",
		16#0f42# => X"18600001",
		16#0f43# => X"ab9c8129",
		16#0f44# => X"a8638112",
		16#0f45# => X"04002639",
		16#0f46# => X"d401e000",
		16#0f47# => X"04001652",
		16#0f48# => X"15000000",
		16#0f49# => X"bc0b0000",
		16#0f4a# => X"0c000344",
		16#0f4b# => X"15000000",
		16#0f4c# => X"0400164d",
		16#0f4d# => X"1a800001",
		16#0f4e# => X"18600001",
		16#0f4f# => X"d4015800",
		16#0f50# => X"0400262e",
		16#0f51# => X"a8637ebc",
		16#0f52# => X"18600001",
		16#0f53# => X"84820000",
		16#0f54# => X"a863819e",
		16#0f55# => X"aa9481b0",
		16#0f56# => X"d4012004",
		16#0f57# => X"04002627",
		16#0f58# => X"d401a000",
		16#0f59# => X"04001640",
		16#0f5a# => X"15000000",
		16#0f5b# => X"bc0b0000",
		16#0f5c# => X"0c000388",
		16#0f5d# => X"15000000",
		16#0f5e# => X"0400163b",
		16#0f5f# => X"1b000001",
		16#0f60# => X"18600001",
		16#0f61# => X"d4015800",
		16#0f62# => X"0400261c",
		16#0f63# => X"a8637ebc",
		16#0f64# => X"18600001",
		16#0f65# => X"ab1881d7",
		16#0f66# => X"a86381c0",
		16#0f67# => X"04002617",
		16#0f68# => X"d401c000",
		16#0f69# => X"04001630",
		16#0f6a# => X"15000000",
		16#0f6b# => X"bc0b0000",
		16#0f6c# => X"0c00031c",
		16#0f6d# => X"15000000",
		16#0f6e# => X"0400162b",
		16#0f6f# => X"15000000",
		16#0f70# => X"18600001",
		16#0f71# => X"d4015800",
		16#0f72# => X"0400260c",
		16#0f73# => X"a8637ebc",
		16#0f74# => X"18600001",
		16#0f75# => X"d401b000",
		16#0f76# => X"04002608",
		16#0f77# => X"a86381dd",
		16#0f78# => X"84a10040",
		16#0f79# => X"a4650001",
		16#0f7a# => X"bc230000",
		16#0f7b# => X"10000285",
		16#0f7c# => X"15000000",
		16#0f7d# => X"84820000",
		16#0f7e# => X"a4650002",
		16#0f7f# => X"bc030000",
		16#0f80# => X"100001ed",
		16#0f81# => X"bc040000",
		16#0f82# => X"100001eb",
		16#0f83# => X"9dc00000",
		16#0f84# => X"00000017",
		16#0f85# => X"9e00004c",
		16#0f86# => X"04001613",
		16#0f87# => X"15000000",
		16#0f88# => X"18600001",
		16#0f89# => X"d4015800",
		16#0f8a# => X"040025f4",
		16#0f8b# => X"a8637ebc",
		16#0f8c# => X"e08e8306",
		16#0f8d# => X"9c610280",
		16#0f8e# => X"e0832000",
		16#0f8f# => X"18600001",
		16#0f90# => X"9484fddc",
		16#0f91# => X"a8638214",
		16#0f92# => X"d4017000",
		16#0f93# => X"9dce0001",
		16#0f94# => X"040025ea",
		16#0f95# => X"d4012004",
		16#0f96# => X"84820000",
		16#0f97# => X"a5ceffff",
		16#0f98# => X"e48e2000",
		16#0f99# => X"0c0001d4",
		16#0f9a# => X"84a10040",
		16#0f9b# => X"040015fe",
		16#0f9c# => X"15000000",
		16#0f9d# => X"bc0b0000",
		16#0f9e# => X"13ffffe8",
		16#0f9f# => X"15000000",
		16#0fa0# => X"040015f9",
		16#0fa1# => X"15000000",
		16#0fa2# => X"040015fd",
		16#0fa3# => X"9c6bffff",
		16#0fa4# => X"03ffffe2",
		16#0fa5# => X"15000000",
		16#0fa6# => X"dc011020",
		16#0fa7# => X"dc011022",
		16#0fa8# => X"9c400066",
		16#0fa9# => X"dc011024",
		16#0faa# => X"84410020",
		16#0fab# => X"e4221800",
		16#0fac# => X"13fffd00",
		16#0fad# => X"98410024",
		16#0fae# => X"bc220000",
		16#0faf# => X"13fffcfd",
		16#0fb0# => X"9c600066",
		16#0fb1# => X"9c403415",
		16#0fb2# => X"dc011824",
		16#0fb3# => X"9c600007",
		16#0fb4# => X"dc011020",
		16#0fb5# => X"0400087e",
		16#0fb6# => X"dc011022",
		16#0fb7# => X"b84b0010",
		16#0fb8# => X"b8420090",
		16#0fb9# => X"bc220000",
		16#0fba# => X"0ffffcf9",
		16#0fbb# => X"15000000",
		16#0fbc# => X"03fffcf9",
		16#0fbd# => X"d4011038",
		16#0fbe# => X"13fffec6",
		16#0fbf# => X"15000000",
		16#0fc0# => X"03fffee7",
		16#0fc1# => X"15000000",
		16#0fc2# => X"03fffd17",
		16#0fc3# => X"d40110d0",
		16#0fc4# => X"03fffcff",
		16#0fc5# => X"d4011084",
		16#0fc6# => X"03fffd6b",
		16#0fc7# => X"d4011200",
		16#0fc8# => X"03fffd53",
		16#0fc9# => X"d40111b4",
		16#0fca# => X"03fffd3b",
		16#0fcb# => X"d4011168",
		16#0fcc# => X"03fffd23",
		16#0fcd# => X"d401111c",
		16#0fce# => X"1000032e",
		16#0fcf# => X"bc0b4eaf",
		16#0fd0# => X"0ffffef5",
		16#0fd1# => X"9c60ffff",
		16#0fd2# => X"040015c7",
		16#0fd3# => X"15000000",
		16#0fd4# => X"bc0b0000",
		16#0fd5# => X"0c000372",
		16#0fd6# => X"15000000",
		16#0fd7# => X"040015c2",
		16#0fd8# => X"15000000",
		16#0fd9# => X"18600001",
		16#0fda# => X"d4015800",
		16#0fdb# => X"040025a3",
		16#0fdc# => X"a8637ebc",
		16#0fdd# => X"18600001",
		16#0fde# => X"04002683",
		16#0fdf# => X"a8637f1c",
		16#0fe0# => X"9c800002",
		16#0fe1# => X"000000e6",
		16#0fe2# => X"d4012018",
		16#0fe3# => X"98a10234",
		16#0fe4# => X"84610038",
		16#0fe5# => X"07fffacd",
		16#0fe6# => X"84810240",
		16#0fe7# => X"84410254",
		16#0fe8# => X"a4620002",
		16#0fe9# => X"bc030000",
		16#0fea# => X"13fffe45",
		16#0feb# => X"d4015a58",
		16#0fec# => X"98a10236",
		16#0fed# => X"98410234",
		16#0fee# => X"b8a50010",
		16#0fef# => X"84610038",
		16#0ff0# => X"84810244",
		16#0ff1# => X"e0a51004",
		16#0ff2# => X"04000509",
		16#0ff3# => X"9cc1025c",
		16#0ff4# => X"84410254",
		16#0ff5# => X"a4420004",
		16#0ff6# => X"bc020000",
		16#0ff7# => X"13fffe3c",
		16#0ff8# => X"98810234",
		16#0ff9# => X"84610038",
		16#0ffa# => X"04000618",
		16#0ffb# => X"84a10248",
		16#0ffc# => X"03fffe38",
		16#0ffd# => X"8441003c",
		16#0ffe# => X"988101e8",
		16#0fff# => X"04000613",
		16#1000# => X"84a101fc",
		16#1001# => X"03fffe27",
		16#1002# => X"84410254",
		16#1003# => X"98a101ea",
		16#1004# => X"984101e8",
		16#1005# => X"b8a50010",
		16#1006# => X"848101f8",
		16#1007# => X"e0a51004",
		16#1008# => X"040004f3",
		16#1009# => X"9cc10210",
		16#100a# => X"03fffe19",
		16#100b# => X"84410208",
		16#100c# => X"98a101e8",
		16#100d# => X"07fffaa5",
		16#100e# => X"848101f4",
		16#100f# => X"84410208",
		16#1010# => X"03fffe0f",
		16#1011# => X"d4015a0c",
		16#1012# => X"9881019c",
		16#1013# => X"040005ff",
		16#1014# => X"84a101b0",
		16#1015# => X"03fffe06",
		16#1016# => X"84410208",
		16#1017# => X"98a1019e",
		16#1018# => X"9841019c",
		16#1019# => X"b8a50010",
		16#101a# => X"848101ac",
		16#101b# => X"e0a51004",
		16#101c# => X"040004df",
		16#101d# => X"9cc101c4",
		16#101e# => X"03fffdf8",
		16#101f# => X"844101bc",
		16#1020# => X"98a1019c",
		16#1021# => X"07fffa91",
		16#1022# => X"848101a8",
		16#1023# => X"844101bc",
		16#1024# => X"03fffdee",
		16#1025# => X"d40159c0",
		16#1026# => X"98810150",
		16#1027# => X"040005eb",
		16#1028# => X"84a10164",
		16#1029# => X"03fffde5",
		16#102a# => X"844101bc",
		16#102b# => X"98a10022",
		16#102c# => X"98410020",
		16#102d# => X"b8a50010",
		16#102e# => X"84610038",
		16#102f# => X"84810030",
		16#1030# => X"e0a51004",
		16#1031# => X"040004ca",
		16#1032# => X"9cc10048",
		16#1033# => X"84410040",
		16#1034# => X"a4420004",
		16#1035# => X"bc020000",
		16#1036# => X"13fffdab",
		16#1037# => X"8441008c",
		16#1038# => X"98810020",
		16#1039# => X"84610038",
		16#103a# => X"040005d8",
		16#103b# => X"84a10034",
		16#103c# => X"8441008c",
		16#103d# => X"a4620001",
		16#103e# => X"bc030000",
		16#103f# => X"13fffda6",
		16#1040# => X"a4620002",
		16#1041# => X"98a1006c",
		16#1042# => X"84610038",
		16#1043# => X"07fffa6f",
		16#1044# => X"84810078",
		16#1045# => X"8441008c",
		16#1046# => X"a4620002",
		16#1047# => X"bc030000",
		16#1048# => X"13fffda0",
		16#1049# => X"d4015890",
		16#104a# => X"98a1006e",
		16#104b# => X"9841006c",
		16#104c# => X"b8a50010",
		16#104d# => X"84610038",
		16#104e# => X"8481007c",
		16#104f# => X"e0a51004",
		16#1050# => X"040004ab",
		16#1051# => X"9cc10094",
		16#1052# => X"8441008c",
		16#1053# => X"a4420004",
		16#1054# => X"bc020000",
		16#1055# => X"13fffd97",
		16#1056# => X"844100d8",
		16#1057# => X"9881006c",
		16#1058# => X"84610038",
		16#1059# => X"040005b9",
		16#105a# => X"84a10080",
		16#105b# => X"844100d8",
		16#105c# => X"a4620001",
		16#105d# => X"bc030000",
		16#105e# => X"13fffd92",
		16#105f# => X"a4620002",
		16#1060# => X"98a100b8",
		16#1061# => X"84610038",
		16#1062# => X"07fffa50",
		16#1063# => X"848100c4",
		16#1064# => X"844100d8",
		16#1065# => X"a4620002",
		16#1066# => X"bc030000",
		16#1067# => X"13fffd8c",
		16#1068# => X"d40158dc",
		16#1069# => X"98a100ba",
		16#106a# => X"984100b8",
		16#106b# => X"b8a50010",
		16#106c# => X"84610038",
		16#106d# => X"848100c8",
		16#106e# => X"e0a51004",
		16#106f# => X"0400048c",
		16#1070# => X"9cc100e0",
		16#1071# => X"844100d8",
		16#1072# => X"a4420004",
		16#1073# => X"bc020000",
		16#1074# => X"13fffd83",
		16#1075# => X"84410124",
		16#1076# => X"988100b8",
		16#1077# => X"84610038",
		16#1078# => X"0400059a",
		16#1079# => X"84a100cc",
		16#107a# => X"84410124",
		16#107b# => X"a4620001",
		16#107c# => X"bc030000",
		16#107d# => X"13fffd7e",
		16#107e# => X"a4620002",
		16#107f# => X"98a10104",
		16#1080# => X"84610038",
		16#1081# => X"07fffa31",
		16#1082# => X"84810110",
		16#1083# => X"84410124",
		16#1084# => X"a4620002",
		16#1085# => X"bc030000",
		16#1086# => X"13fffd78",
		16#1087# => X"d4015928",
		16#1088# => X"98a10106",
		16#1089# => X"98410104",
		16#108a# => X"b8a50010",
		16#108b# => X"84610038",
		16#108c# => X"84810114",
		16#108d# => X"e0a51004",
		16#108e# => X"0400046d",
		16#108f# => X"9cc1012c",
		16#1090# => X"84410124",
		16#1091# => X"a4420004",
		16#1092# => X"bc020000",
		16#1093# => X"13fffd6f",
		16#1094# => X"84410170",
		16#1095# => X"98810104",
		16#1096# => X"84610038",
		16#1097# => X"0400057b",
		16#1098# => X"84a10118",
		16#1099# => X"84410170",
		16#109a# => X"a4620001",
		16#109b# => X"bc030000",
		16#109c# => X"13fffd6a",
		16#109d# => X"a4620002",
		16#109e# => X"98a10150",
		16#109f# => X"84610038",
		16#10a0# => X"07fffa12",
		16#10a1# => X"8481015c",
		16#10a2# => X"84410170",
		16#10a3# => X"a4620002",
		16#10a4# => X"bc030000",
		16#10a5# => X"13fffd64",
		16#10a6# => X"d4015974",
		16#10a7# => X"98a10152",
		16#10a8# => X"98410150",
		16#10a9# => X"b8a50010",
		16#10aa# => X"84610038",
		16#10ab# => X"84810160",
		16#10ac# => X"e0a51004",
		16#10ad# => X"0400044e",
		16#10ae# => X"9cc10178",
		16#10af# => X"03fffd5a",
		16#10b0# => X"84410170",
		16#10b1# => X"98a10020",
		16#10b2# => X"07fffa00",
		16#10b3# => X"8481002c",
		16#10b4# => X"84410040",
		16#10b5# => X"03fffd25",
		16#10b6# => X"d4015844",
		16#10b7# => X"040014e2",
		16#10b8# => X"15000000",
		16#10b9# => X"bc0b0000",
		16#10ba# => X"0c00029f",
		16#10bb# => X"15000000",
		16#10bc# => X"040014dd",
		16#10bd# => X"15000000",
		16#10be# => X"18600001",
		16#10bf# => X"d4015800",
		16#10c0# => X"040024be",
		16#10c1# => X"a8637ebc",
		16#10c2# => X"18600001",
		16#10c3# => X"0400259e",
		16#10c4# => X"a8637f4c",
		16#10c5# => X"9c800003",
		16#10c6# => X"d4012018",
		16#10c7# => X"86420000",
		16#10c8# => X"bc120000",
		16#10c9# => X"13fffdfe",
		16#10ca# => X"18600001",
		16#10cb# => X"e0842000",
		16#10cc# => X"a8638378",
		16#10cd# => X"9e400000",
		16#10ce# => X"e0641800",
		16#10cf# => X"9e00004c",
		16#10d0# => X"d4011810",
		16#10d1# => X"18600001",
		16#10d2# => X"a9d20000",
		16#10d3# => X"a8638384",
		16#10d4# => X"e3c41800",
		16#10d5# => X"18600001",
		16#10d6# => X"a8638390",
		16#10d7# => X"0000000d",
		16#10d8# => X"e3841800",
		16#10d9# => X"9c610280",
		16#10da# => X"e0832000",
		16#10db# => X"9884fde0",
		16#10dc# => X"e2449000",
		16#10dd# => X"9dce0001",
		16#10de# => X"ba520010",
		16#10df# => X"a5ceffff",
		16#10e0# => X"84820000",
		16#10e1# => X"e48e2000",
		16#10e2# => X"0c000062",
		16#10e3# => X"ba520090",
		16#10e4# => X"e0ae8306",
		16#10e5# => X"9c610280",
		16#10e6# => X"e0a32800",
		16#10e7# => X"9c600000",
		16#10e8# => X"8485fdc0",
		16#10e9# => X"a4c40001",
		16#10ea# => X"bc060000",
		16#10eb# => X"10000021",
		16#10ec# => X"dfe51de0",
		16#10ed# => X"84610010",
		16#10ee# => X"94a5fdda",
		16#10ef# => X"97030000",
		16#10f0# => X"e405c000",
		16#10f1# => X"1000001c",
		16#10f2# => X"a4a40002",
		16#10f3# => X"040014a6",
		16#10f4# => X"15000000",
		16#10f5# => X"bc0b0000",
		16#10f6# => X"0c0000fe",
		16#10f7# => X"15000000",
		16#10f8# => X"040014a1",
		16#10f9# => X"e28e8306",
		16#10fa# => X"18600001",
		16#10fb# => X"d4015800",
		16#10fc# => X"04002482",
		16#10fd# => X"a8637ebc",
		16#10fe# => X"9c610280",
		16#10ff# => X"e283a000",
		16#1100# => X"18600001",
		16#1101# => X"9494fdda",
		16#1102# => X"a8637fa3",
		16#1103# => X"d4012004",
		16#1104# => X"d4017000",
		16#1105# => X"04002479",
		16#1106# => X"d401c008",
		16#1107# => X"9cb4fde0",
		16#1108# => X"8494fdc0",
		16#1109# => X"94c50000",
		16#110a# => X"9cc60001",
		16#110b# => X"dc053000",
		16#110c# => X"a4a40002",
		16#110d# => X"bc050000",
		16#110e# => X"10000022",
		16#110f# => X"e0ae8306",
		16#1110# => X"9c610280",
		16#1111# => X"971e0000",
		16#1112# => X"e0a32800",
		16#1113# => X"94a5fddc",
		16#1114# => X"e405c000",
		16#1115# => X"1000001c",
		16#1116# => X"a4840004",
		16#1117# => X"04001482",
		16#1118# => X"15000000",
		16#1119# => X"bc0b0000",
		16#111a# => X"0c0000d4",
		16#111b# => X"15000000",
		16#111c# => X"0400147d",
		16#111d# => X"e28e8306",
		16#111e# => X"18600001",
		16#111f# => X"d4015800",
		16#1120# => X"0400245e",
		16#1121# => X"a8637ebc",
		16#1122# => X"9c610280",
		16#1123# => X"e283a000",
		16#1124# => X"18600001",
		16#1125# => X"9494fddc",
		16#1126# => X"a8637fd2",
		16#1127# => X"d4012004",
		16#1128# => X"d4017000",
		16#1129# => X"04002455",
		16#112a# => X"d401c008",
		16#112b# => X"9cb4fde0",
		16#112c# => X"8494fdc0",
		16#112d# => X"94c50000",
		16#112e# => X"9cc60001",
		16#112f# => X"dc053000",
		16#1130# => X"a4840004",
		16#1131# => X"bc240000",
		16#1132# => X"0fffffa7",
		16#1133# => X"e08e8306",
		16#1134# => X"9c610280",
		16#1135# => X"969c0000",
		16#1136# => X"e0832000",
		16#1137# => X"94a4fdde",
		16#1138# => X"e425a000",
		16#1139# => X"10000019",
		16#113a# => X"15000000",
		16#113b# => X"9884fde0",
		16#113c# => X"e2449000",
		16#113d# => X"9dce0001",
		16#113e# => X"ba520010",
		16#113f# => X"a5ceffff",
		16#1140# => X"84820000",
		16#1141# => X"e48e2000",
		16#1142# => X"13ffffa2",
		16#1143# => X"ba520090",
		16#1144# => X"04000a43",
		16#1145# => X"a652ffff",
		16#1146# => X"04001453",
		16#1147# => X"e24b9000",
		16#1148# => X"ba520010",
		16#1149# => X"bc0b0000",
		16#114a# => X"13fffd85",
		16#114b# => X"ba520090",
		16#114c# => X"0400144d",
		16#114d# => X"15000000",
		16#114e# => X"04001451",
		16#114f# => X"9c6bffff",
		16#1150# => X"03fffd7f",
		16#1151# => X"15000000",
		16#1152# => X"04001447",
		16#1153# => X"15000000",
		16#1154# => X"bc0b0000",
		16#1155# => X"0c0000a5",
		16#1156# => X"15000000",
		16#1157# => X"04001442",
		16#1158# => X"e30e8306",
		16#1159# => X"18600001",
		16#115a# => X"d4015800",
		16#115b# => X"04002423",
		16#115c# => X"a8637ebc",
		16#115d# => X"9c610280",
		16#115e# => X"e303c000",
		16#115f# => X"18600001",
		16#1160# => X"9498fdde",
		16#1161# => X"a8638003",
		16#1162# => X"d4012004",
		16#1163# => X"d4017000",
		16#1164# => X"0400241a",
		16#1165# => X"d401a008",
		16#1166# => X"9cb8fde0",
		16#1167# => X"94850000",
		16#1168# => X"9c840001",
		16#1169# => X"b8840010",
		16#116a# => X"b8840090",
		16#116b# => X"03ffff71",
		16#116c# => X"dc052000",
		16#116d# => X"a4a50004",
		16#116e# => X"bc050000",
		16#116f# => X"1000005a",
		16#1170# => X"9dc00000",
		16#1171# => X"e4247000",
		16#1172# => X"10000019",
		16#1173# => X"9e00004c",
		16#1174# => X"00000022",
		16#1175# => X"bc320000",
		16#1176# => X"04001423",
		16#1177# => X"15000000",
		16#1178# => X"18600001",
		16#1179# => X"d4015800",
		16#117a# => X"04002404",
		16#117b# => X"a8637ebc",
		16#117c# => X"e08e8306",
		16#117d# => X"9c610280",
		16#117e# => X"e0832000",
		16#117f# => X"18600001",
		16#1180# => X"9484fdde",
		16#1181# => X"a8638230",
		16#1182# => X"d4017000",
		16#1183# => X"9dce0001",
		16#1184# => X"040023fa",
		16#1185# => X"d4012004",
		16#1186# => X"84820000",
		16#1187# => X"a5ceffff",
		16#1188# => X"e48e2000",
		16#1189# => X"0c00003f",
		16#118a# => X"15000000",
		16#118b# => X"0400140e",
		16#118c# => X"15000000",
		16#118d# => X"bc0b0000",
		16#118e# => X"13ffffe8",
		16#118f# => X"15000000",
		16#1190# => X"04001409",
		16#1191# => X"15000000",
		16#1192# => X"0400140d",
		16#1193# => X"9c6bffff",
		16#1194# => X"03ffffe2",
		16#1195# => X"15000000",
		16#1196# => X"0c000091",
		16#1197# => X"bdb20000",
		16#1198# => X"10000152",
		16#1199# => X"bd720000",
		16#119a# => X"040013ff",
		16#119b# => X"15000000",
		16#119c# => X"bc0b0000",
		16#119d# => X"0c000192",
		16#119e# => X"15000000",
		16#119f# => X"040013fa",
		16#11a0# => X"15000000",
		16#11a1# => X"18600001",
		16#11a2# => X"d4015800",
		16#11a3# => X"040023db",
		16#11a4# => X"a8637ebc",
		16#11a5# => X"18600001",
		16#11a6# => X"040024bb",
		16#11a7# => X"a86382da",
		16#11a8# => X"04000a01",
		16#11a9# => X"84610028",
		16#11aa# => X"040009ff",
		16#11ab# => X"84610074",
		16#11ac# => X"040009fd",
		16#11ad# => X"846100c0",
		16#11ae# => X"040009fb",
		16#11af# => X"8461010c",
		16#11b0# => X"040009f9",
		16#11b1# => X"84610158",
		16#11b2# => X"040009f7",
		16#11b3# => X"846101a4",
		16#11b4# => X"040009f5",
		16#11b5# => X"846101f0",
		16#11b6# => X"040009f3",
		16#11b7# => X"8461023c",
		16#11b8# => X"04000a81",
		16#11b9# => X"9c610064",
		16#11ba# => X"9c2102ac",
		16#11bb# => X"9d600000",
		16#11bc# => X"8521fffc",
		16#11bd# => X"8441ffd4",
		16#11be# => X"85c1ffd8",
		16#11bf# => X"8601ffdc",
		16#11c0# => X"8641ffe0",
		16#11c1# => X"8681ffe4",
		16#11c2# => X"86c1ffe8",
		16#11c3# => X"8701ffec",
		16#11c4# => X"8741fff0",
		16#11c5# => X"8781fff4",
		16#11c6# => X"44004800",
		16#11c7# => X"87c1fff8",
		16#11c8# => X"9dc00000",
		16#11c9# => X"e4247000",
		16#11ca# => X"10000019",
		16#11cb# => X"9e00004c",
		16#11cc# => X"03ffffca",
		16#11cd# => X"bc320000",
		16#11ce# => X"040013cb",
		16#11cf# => X"15000000",
		16#11d0# => X"18600001",
		16#11d1# => X"d4015800",
		16#11d2# => X"040023ac",
		16#11d3# => X"a8637ebc",
		16#11d4# => X"e08e8306",
		16#11d5# => X"9c610280",
		16#11d6# => X"e0832000",
		16#11d7# => X"18600001",
		16#11d8# => X"9484fdd8",
		16#11d9# => X"a863824c",
		16#11da# => X"d4017000",
		16#11db# => X"9dce0001",
		16#11dc# => X"040023a2",
		16#11dd# => X"d4012004",
		16#11de# => X"84820000",
		16#11df# => X"a5ceffff",
		16#11e0# => X"e48e2000",
		16#11e1# => X"0fffffb5",
		16#11e2# => X"bc320000",
		16#11e3# => X"040013b6",
		16#11e4# => X"15000000",
		16#11e5# => X"bc0b0000",
		16#11e6# => X"13ffffe8",
		16#11e7# => X"15000000",
		16#11e8# => X"040013b1",
		16#11e9# => X"15000000",
		16#11ea# => X"040013b5",
		16#11eb# => X"9c6bffff",
		16#11ec# => X"03ffffe2",
		16#11ed# => X"15000000",
		16#11ee# => X"040013ab",
		16#11ef# => X"15000000",
		16#11f0# => X"040013af",
		16#11f1# => X"9c6bffff",
		16#11f2# => X"03ffff2a",
		16#11f3# => X"15000000",
		16#11f4# => X"040013a5",
		16#11f5# => X"15000000",
		16#11f6# => X"040013a9",
		16#11f7# => X"9c6bffff",
		16#11f8# => X"03ffff00",
		16#11f9# => X"15000000",
		16#11fa# => X"0400139f",
		16#11fb# => X"15000000",
		16#11fc# => X"040013a3",
		16#11fd# => X"9c6bffff",
		16#11fe# => X"03ffff59",
		16#11ff# => X"15000000",
		16#1200# => X"84820000",
		16#1201# => X"bc040000",
		16#1202# => X"13fffd7d",
		16#1203# => X"a4650002",
		16#1204# => X"9dc00000",
		16#1205# => X"00000017",
		16#1206# => X"9e00004c",
		16#1207# => X"04001392",
		16#1208# => X"15000000",
		16#1209# => X"18600001",
		16#120a# => X"d4015800",
		16#120b# => X"04002373",
		16#120c# => X"a8637ebc",
		16#120d# => X"e08e8306",
		16#120e# => X"9c610280",
		16#120f# => X"e0832000",
		16#1210# => X"18600001",
		16#1211# => X"9484fdda",
		16#1212# => X"a86381f8",
		16#1213# => X"d4017000",
		16#1214# => X"9dce0001",
		16#1215# => X"04002369",
		16#1216# => X"d4012004",
		16#1217# => X"84820000",
		16#1218# => X"a5ceffff",
		16#1219# => X"e48e2000",
		16#121a# => X"0ffffd64",
		16#121b# => X"84a10040",
		16#121c# => X"0400137d",
		16#121d# => X"15000000",
		16#121e# => X"bc0b0000",
		16#121f# => X"13ffffe8",
		16#1220# => X"15000000",
		16#1221# => X"04001378",
		16#1222# => X"15000000",
		16#1223# => X"0400137c",
		16#1224# => X"9c6bffff",
		16#1225# => X"03ffffe2",
		16#1226# => X"15000000",
		16#1227# => X"04001372",
		16#1228# => X"15000000",
		16#1229# => X"bc0b0000",
		16#122a# => X"0c000117",
		16#122b# => X"15000000",
		16#122c# => X"0400136d",
		16#122d# => X"15000000",
		16#122e# => X"18600001",
		16#122f# => X"d4015800",
		16#1230# => X"0400234e",
		16#1231# => X"a8637ebc",
		16#1232# => X"18600001",
		16#1233# => X"0400242e",
		16#1234# => X"a8638268",
		16#1235# => X"84610018",
		16#1236# => X"bc230003",
		16#1237# => X"13ffff71",
		16#1238# => X"15000000",
		16#1239# => X"04001360",
		16#123a# => X"15000000",
		16#123b# => X"bc0b0000",
		16#123c# => X"0c000141",
		16#123d# => X"15000000",
		16#123e# => X"0400135b",
		16#123f# => X"15000000",
		16#1240# => X"18600001",
		16#1241# => X"d4015800",
		16#1242# => X"0400233c",
		16#1243# => X"a8637ebc",
		16#1244# => X"84820000",
		16#1245# => X"8461003c",
		16#1246# => X"04001de2",
		16#1247# => X"e0641b06",
		16#1248# => X"d4015810",
		16#1249# => X"d4016014",
		16#124a# => X"0400098f",
		16#124b# => X"a87a0000",
		16#124c# => X"84610010",
		16#124d# => X"84810014",
		16#124e# => X"e0ab0004",
		16#124f# => X"e0cc0004",
		16#1250# => X"04001bbc",
		16#1251# => X"15000000",
		16#1252# => X"18600001",
		16#1253# => X"d4015800",
		16#1254# => X"d4016004",
		16#1255# => X"a86382b1",
		16#1256# => X"d401f008",
		16#1257# => X"04002327",
		16#1258# => X"d401e00c",
		16#1259# => X"04001340",
		16#125a# => X"15000000",
		16#125b# => X"bc0b0000",
		16#125c# => X"0c00011b",
		16#125d# => X"15000000",
		16#125e# => X"0400133b",
		16#125f# => X"15000000",
		16#1260# => X"18600001",
		16#1261# => X"d4015800",
		16#1262# => X"0400231c",
		16#1263# => X"a8637ebc",
		16#1264# => X"18600001",
		16#1265# => X"d401c000",
		16#1266# => X"04002318",
		16#1267# => X"a86382cb",
		16#1268# => X"04001331",
		16#1269# => X"15000000",
		16#126a# => X"bc0b0000",
		16#126b# => X"0c000106",
		16#126c# => X"15000000",
		16#126d# => X"0400132c",
		16#126e# => X"15000000",
		16#126f# => X"18600001",
		16#1270# => X"d4015800",
		16#1271# => X"0400230d",
		16#1272# => X"a8637ebc",
		16#1273# => X"18600001",
		16#1274# => X"84420000",
		16#1275# => X"a86382d1",
		16#1276# => X"d401a004",
		16#1277# => X"04002307",
		16#1278# => X"d4011000",
		16#1279# => X"04001320",
		16#127a# => X"15000000",
		16#127b# => X"bc0b0000",
		16#127c# => X"0c0000ef",
		16#127d# => X"15000000",
		16#127e# => X"0400131b",
		16#127f# => X"15000000",
		16#1280# => X"18600001",
		16#1281# => X"d4015800",
		16#1282# => X"040022fc",
		16#1283# => X"a8637ebc",
		16#1284# => X"0400230e",
		16#1285# => X"9c60000a",
		16#1286# => X"03ffff22",
		16#1287# => X"15000000",
		16#1288# => X"04001311",
		16#1289# => X"15000000",
		16#128a# => X"04001315",
		16#128b# => X"9c6bffff",
		16#128c# => X"03fffce2",
		16#128d# => X"15000000",
		16#128e# => X"0400130b",
		16#128f# => X"15000000",
		16#1290# => X"0400130f",
		16#1291# => X"9c6bffff",
		16#1292# => X"03fffcba",
		16#1293# => X"15000000",
		16#1294# => X"04001305",
		16#1295# => X"15000000",
		16#1296# => X"04001309",
		16#1297# => X"9c6bffff",
		16#1298# => X"03fffca4",
		16#1299# => X"15000000",
		16#129a# => X"040012ff",
		16#129b# => X"15000000",
		16#129c# => X"04001303",
		16#129d# => X"9c6bffff",
		16#129e# => X"03fffc8e",
		16#129f# => X"15000000",
		16#12a0# => X"040012f9",
		16#12a1# => X"15000000",
		16#12a2# => X"040012fd",
		16#12a3# => X"9c6bffff",
		16#12a4# => X"03fffc76",
		16#12a5# => X"15000000",
		16#12a6# => X"040012f3",
		16#12a7# => X"15000000",
		16#12a8# => X"bc0b0000",
		16#12a9# => X"0c00008c",
		16#12aa# => X"15000000",
		16#12ab# => X"040012ee",
		16#12ac# => X"9e520001",
		16#12ad# => X"18600001",
		16#12ae# => X"d4015800",
		16#12af# => X"040022cf",
		16#12b0# => X"a8637ebc",
		16#12b1# => X"18600001",
		16#12b2# => X"ba520010",
		16#12b3# => X"a8638091",
		16#12b4# => X"040023ad",
		16#12b5# => X"ba520090",
		16#12b6# => X"03fffc5f",
		16#12b7# => X"15000000",
		16#12b8# => X"040012e1",
		16#12b9# => X"15000000",
		16#12ba# => X"bc0b0000",
		16#12bb# => X"0c000080",
		16#12bc# => X"15000000",
		16#12bd# => X"040012dc",
		16#12be# => X"15000000",
		16#12bf# => X"18600001",
		16#12c0# => X"d4015800",
		16#12c1# => X"040022bd",
		16#12c2# => X"a8637ebc",
		16#12c3# => X"84820000",
		16#12c4# => X"8461003c",
		16#12c5# => X"04001d63",
		16#12c6# => X"e0641b06",
		16#12c7# => X"d4015810",
		16#12c8# => X"d4016014",
		16#12c9# => X"04000910",
		16#12ca# => X"a87a0000",
		16#12cb# => X"84610010",
		16#12cc# => X"84810014",
		16#12cd# => X"e0ab0004",
		16#12ce# => X"e0cc0004",
		16#12cf# => X"04001b3d",
		16#12d0# => X"15000000",
		16#12d1# => X"18600001",
		16#12d2# => X"d4015800",
		16#12d3# => X"d4016004",
		16#12d4# => X"040022aa",
		16#12d5# => X"a863807a",
		16#12d6# => X"03fffc32",
		16#12d7# => X"15000000",
		16#12d8# => X"040012c1",
		16#12d9# => X"15000000",
		16#12da# => X"040012c5",
		16#12db# => X"9c6bffff",
		16#12dc# => X"03fffc12",
		16#12dd# => X"15000000",
		16#12de# => X"040012bb",
		16#12df# => X"15000000",
		16#12e0# => X"040012bf",
		16#12e1# => X"9c6bffff",
		16#12e2# => X"03fffbfd",
		16#12e3# => X"15000000",
		16#12e4# => X"040012b5",
		16#12e5# => X"15000000",
		16#12e6# => X"040012b9",
		16#12e7# => X"9c6bffff",
		16#12e8# => X"03fffc76",
		16#12e9# => X"15000000",
		16#12ea# => X"13fffebe",
		16#12eb# => X"15000000",
		16#12ec# => X"040012ad",
		16#12ed# => X"15000000",
		16#12ee# => X"bc0b0000",
		16#12ef# => X"0c000076",
		16#12f0# => X"15000000",
		16#12f1# => X"040012a8",
		16#12f2# => X"15000000",
		16#12f3# => X"18600001",
		16#12f4# => X"d4015800",
		16#12f5# => X"04002289",
		16#12f6# => X"a8637ebc",
		16#12f7# => X"18600001",
		16#12f8# => X"04002369",
		16#12f9# => X"a86382ea",
		16#12fa# => X"03fffeae",
		16#12fb# => X"15000000",
		16#12fc# => X"0400129d",
		16#12fd# => X"15000000",
		16#12fe# => X"bc0b0000",
		16#12ff# => X"0c00004e",
		16#1300# => X"15000000",
		16#1301# => X"04001298",
		16#1302# => X"15000000",
		16#1303# => X"18600001",
		16#1304# => X"d4015800",
		16#1305# => X"04002279",
		16#1306# => X"a8637ebc",
		16#1307# => X"18600001",
		16#1308# => X"04002359",
		16#1309# => X"a8637f78",
		16#130a# => X"9c800004",
		16#130b# => X"03fffdbc",
		16#130c# => X"d4012018",
		16#130d# => X"0400128c",
		16#130e# => X"15000000",
		16#130f# => X"bc0b0000",
		16#1310# => X"0c000043",
		16#1311# => X"15000000",
		16#1312# => X"04001287",
		16#1313# => X"15000000",
		16#1314# => X"18600001",
		16#1315# => X"d4015800",
		16#1316# => X"04002268",
		16#1317# => X"a8637ebc",
		16#1318# => X"18600001",
		16#1319# => X"04002348",
		16#131a# => X"a8637ef1",
		16#131b# => X"9c800001",
		16#131c# => X"03fffdab",
		16#131d# => X"d4012018",
		16#131e# => X"0400127b",
		16#131f# => X"15000000",
		16#1320# => X"bc0b0000",
		16#1321# => X"0c00003e",
		16#1322# => X"15000000",
		16#1323# => X"04001276",
		16#1324# => X"15000000",
		16#1325# => X"18600001",
		16#1326# => X"d4015800",
		16#1327# => X"04002257",
		16#1328# => X"a8637ebc",
		16#1329# => X"18600001",
		16#132a# => X"04002337",
		16#132b# => X"a8637ec5",
		16#132c# => X"9c800000",
		16#132d# => X"03fffd9a",
		16#132e# => X"d4012018",
		16#132f# => X"0400126a",
		16#1330# => X"15000000",
		16#1331# => X"0400126e",
		16#1332# => X"9c6bffff",
		16#1333# => X"03fffe6c",
		16#1334# => X"15000000",
		16#1335# => X"04001264",
		16#1336# => X"15000000",
		16#1337# => X"04001268",
		16#1338# => X"9c6bffff",
		16#1339# => X"03ffff72",
		16#133a# => X"15000000",
		16#133b# => X"0400125e",
		16#133c# => X"15000000",
		16#133d# => X"04001262",
		16#133e# => X"9c6bffff",
		16#133f# => X"03ffff7e",
		16#1340# => X"15000000",
		16#1341# => X"04001258",
		16#1342# => X"15000000",
		16#1343# => X"0400125c",
		16#1344# => X"9c6bffff",
		16#1345# => X"03fffee7",
		16#1346# => X"15000000",
		16#1347# => X"04001252",
		16#1348# => X"15000000",
		16#1349# => X"04001256",
		16#134a# => X"9c6bffff",
		16#134b# => X"03fffc8c",
		16#134c# => X"15000000",
		16#134d# => X"0400124c",
		16#134e# => X"15000000",
		16#134f# => X"04001250",
		16#1350# => X"9c6bffff",
		16#1351# => X"03ffffb0",
		16#1352# => X"15000000",
		16#1353# => X"04001246",
		16#1354# => X"15000000",
		16#1355# => X"0400124a",
		16#1356# => X"9c6bffff",
		16#1357# => X"03ffffbb",
		16#1358# => X"15000000",
		16#1359# => X"04001240",
		16#135a# => X"15000000",
		16#135b# => X"04001244",
		16#135c# => X"9c6bffff",
		16#135d# => X"03fffd5f",
		16#135e# => X"15000000",
		16#135f# => X"0400123a",
		16#1360# => X"15000000",
		16#1361# => X"0400123e",
		16#1362# => X"9c6bffff",
		16#1363# => X"03ffffc0",
		16#1364# => X"15000000",
		16#1365# => X"04001234",
		16#1366# => X"15000000",
		16#1367# => X"04001238",
		16#1368# => X"9c6bffff",
		16#1369# => X"03ffff88",
		16#136a# => X"15000000",
		16#136b# => X"0400122e",
		16#136c# => X"15000000",
		16#136d# => X"04001232",
		16#136e# => X"9c6bffff",
		16#136f# => X"03ffff0f",
		16#1370# => X"15000000",
		16#1371# => X"04001228",
		16#1372# => X"15000000",
		16#1373# => X"0400122c",
		16#1374# => X"9c6bffff",
		16#1375# => X"03fffef8",
		16#1376# => X"15000000",
		16#1377# => X"04001222",
		16#1378# => X"15000000",
		16#1379# => X"04001226",
		16#137a# => X"9c6bffff",
		16#137b# => X"03fffee3",
		16#137c# => X"15000000",
		16#137d# => X"0400121c",
		16#137e# => X"15000000",
		16#137f# => X"04001220",
		16#1380# => X"9c6bffff",
		16#1381# => X"03fffebd",
		16#1382# => X"15000000",
		16#1383# => X"b8e70010",
		16#1384# => X"d7e117d4",
		16#1385# => X"d7e187dc",
		16#1386# => X"d7e1d7f0",
		16#1387# => X"d7e1e7f4",
		16#1388# => X"d7e1f7f8",
		16#1389# => X"d7e14ffc",
		16#138a# => X"d7e177d8",
		16#138b# => X"d7e197e0",
		16#138c# => X"d7e1a7e4",
		16#138d# => X"d7e1b7e8",
		16#138e# => X"d7e1c7ec",
		16#138f# => X"a8430000",
		16#1390# => X"9c21ffd4",
		16#1391# => X"ab840000",
		16#1392# => X"abc50000",
		16#1393# => X"ab460000",
		16#1394# => X"bc030000",
		16#1395# => X"10000147",
		16#1396# => X"ba070090",
		16#1397# => X"a690ffff",
		16#1398# => X"e1c31800",
		16#1399# => X"aac50000",
		16#139a# => X"a9650000",
		16#139b# => X"9cc00000",
		16#139c# => X"a86b0000",
		16#139d# => X"9ce00000",
		16#139e# => X"95030000",
		16#139f# => X"e1144000",
		16#13a0# => X"9ce70001",
		16#13a1# => X"dc034000",
		16#13a2# => X"e4423800",
		16#13a3# => X"13fffffb",
		16#13a4# => X"9c630002",
		16#13a5# => X"9cc60001",
		16#13a6# => X"e4423000",
		16#13a7# => X"13fffff5",
		16#13a8# => X"e16b7000",
		16#13a9# => X"ba420002",
		16#13aa# => X"ab1c0000",
		16#13ab# => X"a9bc0000",
		16#13ac# => X"a99e0000",
		16#13ad# => X"9cc00000",
		16#13ae# => X"a90d0000",
		16#13af# => X"a8ec0000",
		16#13b0# => X"9c600000",
		16#13b1# => X"99670000",
		16#13b2# => X"e1705b06",
		16#13b3# => X"9c630001",
		16#13b4# => X"d4085800",
		16#13b5# => X"9ce70002",
		16#13b6# => X"e4421800",
		16#13b7# => X"13fffffa",
		16#13b8# => X"9d080004",
		16#13b9# => X"9cc60001",
		16#13ba# => X"e18c7000",
		16#13bb# => X"e4a23000",
		16#13bc# => X"0ffffff2",
		16#13bd# => X"e1ad9000",
		16#13be# => X"9ee00000",
		16#13bf# => X"9c60f000",
		16#13c0# => X"a8dc0000",
		16#13c1# => X"e2101804",
		16#13c2# => X"a8f70000",
		16#13c3# => X"a8770000",
		16#13c4# => X"a9b70000",
		16#13c5# => X"a9660000",
		16#13c6# => X"aa270000",
		16#13c7# => X"9d000000",
		16#13c8# => X"a583ffff",
		16#13c9# => X"84eb0000",
		16#13ca# => X"9e6c000a",
		16#13cb# => X"e5478800",
		16#13cc# => X"ba730010",
		16#13cd# => X"9d080001",
		16#13ce# => X"e06d3800",
		16#13cf# => X"9de00001",
		16#13d0# => X"aa270000",
		16#13d1# => X"10000003",
		16#13d2# => X"ba730090",
		16#13d3# => X"9de00000",
		16#13d4# => X"e18c7800",
		16#13d5# => X"a9a30000",
		16#13d6# => X"b98c0010",
		16#13d7# => X"e5701800",
		16#13d8# => X"9d6b0004",
		16#13d9# => X"10000004",
		16#13da# => X"b98c0090",
		16#13db# => X"9da00000",
		16#13dc# => X"e5701800",
		16#13dd# => X"10000003",
		16#13de# => X"e4424000",
		16#13df# => X"a9930000",
		16#13e0# => X"13ffffe8",
		16#13e1# => X"a86c0000",
		16#13e2# => X"9ef70001",
		16#13e3# => X"e4a2b800",
		16#13e4# => X"0fffffe1",
		16#13e5# => X"e0c69000",
		16#13e6# => X"9c800000",
		16#13e7# => X"040006ec",
		16#13e8# => X"a86c0000",
		16#13e9# => X"aa7e0000",
		16#13ea# => X"a88b0000",
		16#13eb# => X"aa3c0000",
		16#13ec# => X"9cc00000",
		16#13ed# => X"9d800000",
		16#13ee# => X"a91a0000",
		16#13ef# => X"d4116000",
		16#13f0# => X"a8f30000",
		16#13f1# => X"a86c0000",
		16#13f2# => X"99e80000",
		16#13f3# => X"99a70000",
		16#13f4# => X"e1af6b06",
		16#13f5# => X"9c630001",
		16#13f6# => X"e18c6800",
		16#13f7# => X"9ce70002",
		16#13f8# => X"e4421800",
		16#13f9# => X"13fffff9",
		16#13fa# => X"9d080002",
		16#13fb# => X"d4116000",
		16#13fc# => X"9cc60001",
		16#13fd# => X"9e310004",
		16#13fe# => X"e4423000",
		16#13ff# => X"13ffffee",
		16#1400# => X"e2737000",
		16#1401# => X"9ee00000",
		16#1402# => X"a8dc0000",
		16#1403# => X"a8770000",
		16#1404# => X"a8f70000",
		16#1405# => X"a9f70000",
		16#1406# => X"a9860000",
		16#1407# => X"aa670000",
		16#1408# => X"9d000000",
		16#1409# => X"a5a3ffff",
		16#140a# => X"84ec0000",
		16#140b# => X"9ead000a",
		16#140c# => X"e5479800",
		16#140d# => X"bab50010",
		16#140e# => X"9d080001",
		16#140f# => X"e06f3800",
		16#1410# => X"9e200001",
		16#1411# => X"aa670000",
		16#1412# => X"10000003",
		16#1413# => X"bab50090",
		16#1414# => X"9e200000",
		16#1415# => X"e1ad8800",
		16#1416# => X"a9e30000",
		16#1417# => X"b9ad0010",
		16#1418# => X"e5701800",
		16#1419# => X"9d8c0004",
		16#141a# => X"10000004",
		16#141b# => X"b9ad0090",
		16#141c# => X"9de00000",
		16#141d# => X"e5701800",
		16#141e# => X"10000003",
		16#141f# => X"e4424000",
		16#1420# => X"a9b50000",
		16#1421# => X"13ffffe8",
		16#1422# => X"a86d0000",
		16#1423# => X"9ef70001",
		16#1424# => X"e4a2b800",
		16#1425# => X"0fffffe1",
		16#1426# => X"e0c69000",
		16#1427# => X"040006ac",
		16#1428# => X"a86d0000",
		16#1429# => X"ab7c0000",
		16#142a# => X"a88b0000",
		16#142b# => X"aafe0000",
		16#142c# => X"9cc00000",
		16#142d# => X"aaba0000",
		16#142e# => X"aa3b0000",
		16#142f# => X"9e600000",
		16#1430# => X"9d800000",
		16#1431# => X"a9150000",
		16#1432# => X"d4116000",
		16#1433# => X"a8f70000",
		16#1434# => X"a86c0000",
		16#1435# => X"99e80000",
		16#1436# => X"99a70000",
		16#1437# => X"e1af6b06",
		16#1438# => X"9c630001",
		16#1439# => X"e18c6800",
		16#143a# => X"9ce70002",
		16#143b# => X"e4421800",
		16#143c# => X"13fffff9",
		16#143d# => X"e1087000",
		16#143e# => X"d4116000",
		16#143f# => X"9e730001",
		16#1440# => X"9e310004",
		16#1441# => X"e4429800",
		16#1442# => X"13ffffee",
		16#1443# => X"9eb50002",
		16#1444# => X"9cc60001",
		16#1445# => X"e2f77000",
		16#1446# => X"e4423000",
		16#1447# => X"13ffffe6",
		16#1448# => X"e37b9000",
		16#1449# => X"9ee00000",
		16#144a# => X"a8dc0000",
		16#144b# => X"a8770000",
		16#144c# => X"a8f70000",
		16#144d# => X"a9f70000",
		16#144e# => X"a9860000",
		16#144f# => X"aa670000",
		16#1450# => X"9d000000",
		16#1451# => X"a5a3ffff",
		16#1452# => X"84ec0000",
		16#1453# => X"9ead000a",
		16#1454# => X"e5479800",
		16#1455# => X"bab50010",
		16#1456# => X"9d080001",
		16#1457# => X"e06f3800",
		16#1458# => X"9e200001",
		16#1459# => X"aa670000",
		16#145a# => X"10000003",
		16#145b# => X"bab50090",
		16#145c# => X"9e200000",
		16#145d# => X"e1ad8800",
		16#145e# => X"a9e30000",
		16#145f# => X"b9ad0010",
		16#1460# => X"e5701800",
		16#1461# => X"9d8c0004",
		16#1462# => X"10000004",
		16#1463# => X"b9ad0090",
		16#1464# => X"9de00000",
		16#1465# => X"e5701800",
		16#1466# => X"10000003",
		16#1467# => X"e4424000",
		16#1468# => X"a9b50000",
		16#1469# => X"13ffffe8",
		16#146a# => X"a86d0000",
		16#146b# => X"9ef70001",
		16#146c# => X"e4a2b800",
		16#146d# => X"0fffffe1",
		16#146e# => X"e0c69000",
		16#146f# => X"04000664",
		16#1470# => X"a86d0000",
		16#1471# => X"ab3c0000",
		16#1472# => X"a88b0000",
		16#1473# => X"aabe0000",
		16#1474# => X"9ee00000",
		16#1475# => X"aa7a0000",
		16#1476# => X"a9f90000",
		16#1477# => X"9e200000",
		16#1478# => X"9d000000",
		16#1479# => X"a8f30000",
		16#147a# => X"d40f4000",
		16#147b# => X"a8b50000",
		16#147c# => X"a8680000",
		16#147d# => X"99a70000",
		16#147e# => X"99850000",
		16#147f# => X"e18d6306",
		16#1480# => X"b9ac0085",
		16#1481# => X"b98c0082",
		16#1482# => X"9c630001",
		16#1483# => X"a5ad007f",
		16#1484# => X"a58c000f",
		16#1485# => X"9ca50002",
		16#1486# => X"e18d6306",
		16#1487# => X"e0e77000",
		16#1488# => X"e4421800",
		16#1489# => X"13fffff4",
		16#148a# => X"e1086000",
		16#148b# => X"d40f4000",
		16#148c# => X"9e310001",
		16#148d# => X"9def0004",
		16#148e# => X"e4428800",
		16#148f# => X"13ffffe9",
		16#1490# => X"9e730002",
		16#1491# => X"9ef70001",
		16#1492# => X"e2b57000",
		16#1493# => X"e442b800",
		16#1494# => X"13ffffe1",
		16#1495# => X"e3399000",
		16#1496# => X"9e600000",
		16#1497# => X"a8730000",
		16#1498# => X"a8b30000",
		16#1499# => X"a9930000",
		16#149a# => X"a8f80000",
		16#149b# => X"a9e50000",
		16#149c# => X"9cc00000",
		16#149d# => X"a503ffff",
		16#149e# => X"84a70000",
		16#149f# => X"9e28000a",
		16#14a0# => X"e5457800",
		16#14a1# => X"ba310010",
		16#14a2# => X"9cc60001",
		16#14a3# => X"e06c2800",
		16#14a4# => X"9da00001",
		16#14a5# => X"a9e50000",
		16#14a6# => X"10000003",
		16#14a7# => X"ba310090",
		16#14a8# => X"9da00000",
		16#14a9# => X"e1086800",
		16#14aa# => X"a9830000",
		16#14ab# => X"b9080010",
		16#14ac# => X"e5701800",
		16#14ad# => X"9ce70004",
		16#14ae# => X"10000004",
		16#14af# => X"b9080090",
		16#14b0# => X"9d800000",
		16#14b1# => X"e5701800",
		16#14b2# => X"10000003",
		16#14b3# => X"e4423000",
		16#14b4# => X"a9110000",
		16#14b5# => X"13ffffe8",
		16#14b6# => X"a8680000",
		16#14b7# => X"9e730001",
		16#14b8# => X"e4a29800",
		16#14b9# => X"0fffffe1",
		16#14ba# => X"e3189000",
		16#14bb# => X"04000618",
		16#14bc# => X"a8680000",
		16#14bd# => X"e0c0a002",
		16#14be# => X"9ce00000",
		16#14bf# => X"a4c6ffff",
		16#14c0# => X"a8760000",
		16#14c1# => X"9c800000",
		16#14c2# => X"94a30000",
		16#14c3# => X"e0a62800",
		16#14c4# => X"9c840001",
		16#14c5# => X"dc032800",
		16#14c6# => X"e4422000",
		16#14c7# => X"13fffffb",
		16#14c8# => X"9c630002",
		16#14c9# => X"9ce70001",
		16#14ca# => X"e4a23800",
		16#14cb# => X"0ffffff5",
		16#14cc# => X"e2d67000",
		16#14cd# => X"9c21002c",
		16#14ce# => X"b96b0010",
		16#14cf# => X"8521fffc",
		16#14d0# => X"8441ffd4",
		16#14d1# => X"b96b0090",
		16#14d2# => X"85c1ffd8",
		16#14d3# => X"8601ffdc",
		16#14d4# => X"8641ffe0",
		16#14d5# => X"8681ffe4",
		16#14d6# => X"86c1ffe8",
		16#14d7# => X"8701ffec",
		16#14d8# => X"8741fff0",
		16#14d9# => X"8781fff4",
		16#14da# => X"44004800",
		16#14db# => X"87c1fff8",
		16#14dc# => X"040005f7",
		16#14dd# => X"a8830000",
		16#14de# => X"a8620000",
		16#14df# => X"040005f4",
		16#14e0# => X"a88b0000",
		16#14e1# => X"a8620000",
		16#14e2# => X"040005f1",
		16#14e3# => X"a88b0000",
		16#14e4# => X"a8620000",
		16#14e5# => X"040005ee",
		16#14e6# => X"a88b0000",
		16#14e7# => X"03ffffe7",
		16#14e8# => X"9c21002c",
		16#14e9# => X"b8e40010",
		16#14ea# => X"a8c30000",
		16#14eb# => X"d7e14ffc",
		16#14ec# => X"b8e70090",
		16#14ed# => X"d7e117f8",
		16#14ee# => X"8486000c",
		16#14ef# => X"a445ffff",
		16#14f0# => X"9c21fff8",
		16#14f1# => X"84630000",
		16#14f2# => X"84a60004",
		16#14f3# => X"07fffe90",
		16#14f4# => X"84c60008",
		16#14f5# => X"9c210008",
		16#14f6# => X"a8820000",
		16#14f7# => X"a86b0000",
		16#14f8# => X"8521fffc",
		16#14f9# => X"000005da",
		16#14fa# => X"8441fff8",
		16#14fb# => X"d7e117fc",
		16#14fc# => X"bc050000",
		16#14fd# => X"0c000003",
		16#14fe# => X"9c21fffc",
		16#14ff# => X"9ca00001",
		16#1500# => X"bc030000",
		16#1501# => X"0c000005",
		16#1502# => X"9d600000",
		16#1503# => X"0000003b",
		16#1504# => X"9c84ffff",
		16#1505# => X"a9670000",
		16#1506# => X"9ceb0001",
		16#1507# => X"e1073b06",
		16#1508# => X"b9080003",
		16#1509# => X"e4434000",
		16#150a# => X"13fffffb",
		16#150b# => X"e32b5b06",
		16#150c# => X"9c84ffff",
		16#150d# => X"9c40fffc",
		16#150e# => X"e339c800",
		16#150f# => X"e2641003",
		16#1510# => X"bc2b0000",
		16#1511# => X"9e730004",
		16#1512# => X"0c000020",
		16#1513# => X"e2b3c800",
		16#1514# => X"9de00000",
		16#1515# => X"e2eb5800",
		16#1516# => X"aa2f0000",
		16#1517# => X"9c600001",
		16#1518# => X"e1157800",
		16#1519# => X"e0f37800",
		16#151a# => X"9c800000",
		16#151b# => X"e0a51b06",
		16#151c# => X"b985009f",
		16#151d# => X"a5a3ffff",
		16#151e# => X"9c840001",
		16#151f# => X"b98c0050",
		16#1520# => X"9c630001",
		16#1521# => X"e4845800",
		16#1522# => X"e0a56000",
		16#1523# => X"a4a5ffff",
		16#1524# => X"e0a56002",
		16#1525# => X"e18d2800",
		16#1526# => X"a58cffff",
		16#1527# => X"e1ac6800",
		16#1528# => X"dc086000",
		16#1529# => X"a5ad00ff",
		16#152a# => X"9d080002",
		16#152b# => X"dc076800",
		16#152c# => X"13ffffef",
		16#152d# => X"9ce70002",
		16#152e# => X"9e310001",
		16#152f# => X"e4715800",
		16#1530# => X"0fffffe8",
		16#1531# => X"e1efb800",
		16#1532# => X"e075c800",
		16#1533# => X"9c40fffc",
		16#1534# => X"9c63ffff",
		16#1535# => X"9c210004",
		16#1536# => X"e0631003",
		16#1537# => X"d4069804",
		16#1538# => X"9c630004",
		16#1539# => X"d406a808",
		16#153a# => X"d4065800",
		16#153b# => X"d406180c",
		16#153c# => X"44004800",
		16#153d# => X"8441fffc",
		16#153e# => X"9c40fffc",
		16#153f# => X"9f200002",
		16#1540# => X"e2a41003",
		16#1541# => X"9d60ffff",
		16#1542# => X"9e750004",
		16#1543# => X"03ffffd1",
		16#1544# => X"9eb50006",
		16#1545# => X"b8a50010",
		16#1546# => X"a9630000",
		16#1547# => X"bc030000",
		16#1548# => X"10000027",
		16#1549# => X"ba250090",
		16#154a# => X"9ea00000",
		16#154b# => X"bae30002",
		16#154c# => X"a9750000",
		16#154d# => X"a9f50000",
		16#154e# => X"a9950000",
		16#154f# => X"a9040000",
		16#1550# => X"9ce00000",
		16#1551# => X"a56bffff",
		16#1552# => X"84c80000",
		16#1553# => X"9e6b000a",
		16#1554# => X"9ce70001",
		16#1555# => X"ba730010",
		16#1556# => X"e0ac3000",
		16#1557# => X"9da00001",
		16#1558# => X"e5467800",
		16#1559# => X"10000003",
		16#155a# => X"ba730090",
		16#155b# => X"9da00000",
		16#155c# => X"e16b6800",
		16#155d# => X"a9850000",
		16#155e# => X"b96b0010",
		16#155f# => X"e5a58800",
		16#1560# => X"9d080004",
		16#1561# => X"a9e60000",
		16#1562# => X"10000004",
		16#1563# => X"b96b0090",
		16#1564# => X"9d800000",
		16#1565# => X"e5a58800",
		16#1566# => X"10000003",
		16#1567# => X"e4433800",
		16#1568# => X"a9730000",
		16#1569# => X"13ffffe8",
		16#156a# => X"15000000",
		16#156b# => X"9eb50001",
		16#156c# => X"e4a3a800",
		16#156d# => X"0fffffe2",
		16#156e# => X"e084b800",
		16#156f# => X"44004800",
		16#1570# => X"15000000",
		16#1571# => X"b8c60010",
		16#1572# => X"bc030000",
		16#1573# => X"10000015",
		16#1574# => X"b9860090",
		16#1575# => X"b9e30002",
		16#1576# => X"e2231800",
		16#1577# => X"9da00000",
		16#1578# => X"a9040000",
		16#1579# => X"a8e50000",
		16#157a# => X"9cc00000",
		16#157b# => X"99670000",
		16#157c# => X"e16c5b06",
		16#157d# => X"9cc60001",
		16#157e# => X"d4085800",
		16#157f# => X"9ce70002",
		16#1580# => X"e4433000",
		16#1581# => X"13fffffa",
		16#1582# => X"9d080004",
		16#1583# => X"9dad0001",
		16#1584# => X"e0a58800",
		16#1585# => X"e4a36800",
		16#1586# => X"0ffffff2",
		16#1587# => X"e0847800",
		16#1588# => X"44004800",
		16#1589# => X"15000000",
		16#158a# => X"b8a50010",
		16#158b# => X"bc030000",
		16#158c# => X"10000012",
		16#158d# => X"b8a50090",
		16#158e# => X"a505ffff",
		16#158f# => X"e1831800",
		16#1590# => X"9d600000",
		16#1591# => X"a8a40000",
		16#1592# => X"9cc00000",
		16#1593# => X"94e50000",
		16#1594# => X"e0e83800",
		16#1595# => X"9cc60001",
		16#1596# => X"dc053800",
		16#1597# => X"e4433000",
		16#1598# => X"13fffffb",
		16#1599# => X"9ca50002",
		16#159a# => X"9d6b0001",
		16#159b# => X"e4a35800",
		16#159c# => X"0ffffff5",
		16#159d# => X"e0846000",
		16#159e# => X"44004800",
		16#159f# => X"15000000",
		16#15a0# => X"d7e117fc",
		16#15a1# => X"bc030000",
		16#15a2# => X"10000018",
		16#15a3# => X"9c21fffc",
		16#15a4# => X"e2631800",
		16#15a5# => X"9e200000",
		16#15a6# => X"9d800000",
		16#15a7# => X"a9660000",
		16#15a8# => X"d4046000",
		16#15a9# => X"a9050000",
		16#15aa# => X"a8ec0000",
		16#15ab# => X"99eb0000",
		16#15ac# => X"99a80000",
		16#15ad# => X"e1af6b06",
		16#15ae# => X"9ce70001",
		16#15af# => X"e18c6800",
		16#15b0# => X"9d080002",
		16#15b1# => X"e4433800",
		16#15b2# => X"13fffff9",
		16#15b3# => X"9d6b0002",
		16#15b4# => X"d4046000",
		16#15b5# => X"9e310001",
		16#15b6# => X"9c840004",
		16#15b7# => X"e4438800",
		16#15b8# => X"13ffffee",
		16#15b9# => X"e0a59800",
		16#15ba# => X"9c210004",
		16#15bb# => X"44004800",
		16#15bc# => X"8441fffc",
		16#15bd# => X"d7e117fc",
		16#15be# => X"bc030000",
		16#15bf# => X"10000023",
		16#15c0# => X"9c21fffc",
		16#15c1# => X"bb630002",
		16#15c2# => X"e1a31800",
		16#15c3# => X"aaa50000",
		16#15c4# => X"ab240000",
		16#15c5# => X"9ee00000",
		16#15c6# => X"aa660000",
		16#15c7# => X"a9f90000",
		16#15c8# => X"9e200000",
		16#15c9# => X"9d000000",
		16#15ca# => X"a8f30000",
		16#15cb# => X"d40f4000",
		16#15cc# => X"a8b50000",
		16#15cd# => X"a8880000",
		16#15ce# => X"99870000",
		16#15cf# => X"99650000",
		16#15d0# => X"e16c5b06",
		16#15d1# => X"9c840001",
		16#15d2# => X"e1085800",
		16#15d3# => X"9ca50002",
		16#15d4# => X"e4432000",
		16#15d5# => X"13fffff9",
		16#15d6# => X"e0e76800",
		16#15d7# => X"d40f4000",
		16#15d8# => X"9e310001",
		16#15d9# => X"9def0004",
		16#15da# => X"e4438800",
		16#15db# => X"13ffffee",
		16#15dc# => X"9e730002",
		16#15dd# => X"9ef70001",
		16#15de# => X"e2b56800",
		16#15df# => X"e4a3b800",
		16#15e0# => X"0fffffe6",
		16#15e1# => X"e339d800",
		16#15e2# => X"9c210004",
		16#15e3# => X"44004800",
		16#15e4# => X"8441fffc",
		16#15e5# => X"d7e117fc",
		16#15e6# => X"bc030000",
		16#15e7# => X"10000028",
		16#15e8# => X"9c21fffc",
		16#15e9# => X"bb630002",
		16#15ea# => X"e1a31800",
		16#15eb# => X"aaa50000",
		16#15ec# => X"ab240000",
		16#15ed# => X"9ee00000",
		16#15ee# => X"aa660000",
		16#15ef# => X"a9f90000",
		16#15f0# => X"9e200000",
		16#15f1# => X"9d000000",
		16#15f2# => X"a8f30000",
		16#15f3# => X"d40f4000",
		16#15f4# => X"a8b50000",
		16#15f5# => X"a8880000",
		16#15f6# => X"99870000",
		16#15f7# => X"99650000",
		16#15f8# => X"e16c5b06",
		16#15f9# => X"b98b0085",
		16#15fa# => X"b96b0082",
		16#15fb# => X"9c840001",
		16#15fc# => X"a58c007f",
		16#15fd# => X"a56b000f",
		16#15fe# => X"9ca50002",
		16#15ff# => X"e16c5b06",
		16#1600# => X"e0e76800",
		16#1601# => X"e4432000",
		16#1602# => X"13fffff4",
		16#1603# => X"e1085800",
		16#1604# => X"d40f4000",
		16#1605# => X"9e310001",
		16#1606# => X"9def0004",
		16#1607# => X"e4438800",
		16#1608# => X"13ffffe9",
		16#1609# => X"9e730002",
		16#160a# => X"9ef70001",
		16#160b# => X"e2b56800",
		16#160c# => X"e4a3b800",
		16#160d# => X"0fffffe1",
		16#160e# => X"e339d800",
		16#160f# => X"9c210004",
		16#1610# => X"44004800",
		16#1611# => X"8441fffc",
		16#1612# => X"b8840010",
		16#1613# => X"9ce00000",
		16#1614# => X"d7e117fc",
		16#1615# => X"baa40090",
		16#1616# => X"9c21fffc",
		16#1617# => X"9f63ffff",
		16#1618# => X"a9870000",
		16#1619# => X"a9070000",
		16#161a# => X"e3286000",
		16#161b# => X"9ef90001",
		16#161c# => X"e45bb800",
		16#161d# => X"0c000056",
		16#161e# => X"e4a34000",
		16#161f# => X"bc0c0000",
		16#1620# => X"1000003f",
		16#1621# => X"15000000",
		16#1622# => X"ba6c0042",
		16#1623# => X"b8930002",
		16#1624# => X"e1602002",
		16#1625# => X"e16b2004",
		16#1626# => X"ad6bffff",
		16#1627# => X"b96b005f",
		16#1628# => X"bc2b0000",
		16#1629# => X"1000009a",
		16#162a# => X"e1e54000",
		16#162b# => X"bc4c0003",
		16#162c# => X"10000003",
		16#162d# => X"9cc00001",
		16#162e# => X"a8cb0000",
		16#162f# => X"e16f3804",
		16#1630# => X"9fa70004",
		16#1631# => X"a56b0003",
		16#1632# => X"9da00001",
		16#1633# => X"e2205802",
		16#1634# => X"e44fe800",
		16#1635# => X"e1715804",
		16#1636# => X"ad6bffff",
		16#1637# => X"b96b005f",
		16#1638# => X"10000003",
		16#1639# => X"e0c65803",
		16#163a# => X"9da00000",
		16#163b# => X"9e2f0004",
		16#163c# => X"e4478800",
		16#163d# => X"10000003",
		16#163e# => X"9d600001",
		16#163f# => X"9d600000",
		16#1640# => X"e16d5804",
		16#1641# => X"e0c65803",
		16#1642# => X"acc60001",
		16#1643# => X"bc260000",
		16#1644# => X"1000007f",
		16#1645# => X"15000000",
		16#1646# => X"a9660000",
		16#1647# => X"e1a73000",
		16#1648# => X"e22f3000",
		16#1649# => X"85ad0000",
		16#164a# => X"9d6b0001",
		16#164b# => X"d4116800",
		16#164c# => X"e4535800",
		16#164d# => X"13fffffa",
		16#164e# => X"9cc60004",
		16#164f# => X"e40c2000",
		16#1650# => X"1000000b",
		16#1651# => X"15000000",
		16#1652# => X"e1044000",
		16#1653# => X"e1054000",
		16#1654# => X"e0c72000",
		16#1655# => X"9c840001",
		16#1656# => X"8cc60000",
		16#1657# => X"d8083000",
		16#1658# => X"e44c2000",
		16#1659# => X"13fffffb",
		16#165a# => X"9d080001",
		16#165b# => X"e325c800",
		16#165c# => X"9c40002c",
		16#165d# => X"a9170000",
		16#165e# => X"d8191000",
		16#165f# => X"9eb50001",
		16#1660# => X"b8d50010",
		16#1661# => X"baa60090",
		16#1662# => X"a4950007",
		16#1663# => X"9c84fffd",
		16#1664# => X"bc440004",
		16#1665# => X"0c00003e",
		16#1666# => X"18400001",
		16#1667# => X"b8860051",
		16#1668# => X"9d800004",
		16#1669# => X"18400001",
		16#166a# => X"a484000c",
		16#166b# => X"a84283d0",
		16#166c# => X"e3286000",
		16#166d# => X"e0841000",
		16#166e# => X"9ef90001",
		16#166f# => X"e45bb800",
		16#1670# => X"13ffffaf",
		16#1671# => X"84e40000",
		16#1672# => X"e4a34000",
		16#1673# => X"1000002d",
		16#1674# => X"e1634002",
		16#1675# => X"e0e54000",
		16#1676# => X"e0c03802",
		16#1677# => X"a4c60003",
		16#1678# => X"e4a65800",
		16#1679# => X"0c000048",
		16#167a# => X"a9a70000",
		16#167b# => X"bc060000",
		16#167c# => X"1000000e",
		16#167d# => X"9c800000",
		16#167e# => X"00000004",
		16#167f# => X"9c400000",
		16#1680# => X"e0e54000",
		16#1681# => X"9c400000",
		16#1682# => X"9c840001",
		16#1683# => X"d8071000",
		16#1684# => X"e4843000",
		16#1685# => X"13fffffb",
		16#1686# => X"9d080001",
		16#1687# => X"e40b3000",
		16#1688# => X"10000018",
		16#1689# => X"15000000",
		16#168a# => X"e16b3002",
		16#168b# => X"b8eb0042",
		16#168c# => X"b9870002",
		16#168d# => X"bc0c0000",
		16#168e# => X"1000000c",
		16#168f# => X"9c800000",
		16#1690# => X"e0cd3000",
		16#1691# => X"9c400000",
		16#1692# => X"9c840001",
		16#1693# => X"d4061000",
		16#1694# => X"e4843800",
		16#1695# => X"13fffffd",
		16#1696# => X"9cc60004",
		16#1697# => X"e40b6000",
		16#1698# => X"10000008",
		16#1699# => X"e1086000",
		16#169a# => X"e0854000",
		16#169b# => X"9c400000",
		16#169c# => X"9d080001",
		16#169d# => X"e4434000",
		16#169e# => X"13fffffc",
		16#169f# => X"d8041000",
		16#16a0# => X"9c210004",
		16#16a1# => X"44004800",
		16#16a2# => X"8441fffc",
		16#16a3# => X"b8840002",
		16#16a4# => X"a842839c",
		16#16a5# => X"e0841000",
		16#16a6# => X"84840000",
		16#16a7# => X"44002000",
		16#16a8# => X"15000000",
		16#16a9# => X"b8950041",
		16#16aa# => X"18400001",
		16#16ab# => X"9d800008",
		16#16ac# => X"a484000c",
		16#16ad# => X"a84283e0",
		16#16ae# => X"e0841000",
		16#16af# => X"03ffff6b",
		16#16b0# => X"84e40000",
		16#16b1# => X"b8950041",
		16#16b2# => X"18400001",
		16#16b3# => X"9d800008",
		16#16b4# => X"a484000c",
		16#16b5# => X"a84283f0",
		16#16b6# => X"e0841000",
		16#16b7# => X"03ffff63",
		16#16b8# => X"84e40000",
		16#16b9# => X"b8950041",
		16#16ba# => X"18400001",
		16#16bb# => X"9d800008",
		16#16bc# => X"a484000c",
		16#16bd# => X"a8428400",
		16#16be# => X"e0841000",
		16#16bf# => X"03ffff5b",
		16#16c0# => X"84e40000",
		16#16c1# => X"03ffffba",
		16#16c2# => X"a8cb0000",
		16#16c3# => X"03ffff8f",
		16#16c4# => X"9c800000",
		16#16c5# => X"d7e117fc",
		16#16c6# => X"84c30000",
		16#16c7# => X"8ca60000",
		16#16c8# => X"e1602802",
		16#16c9# => X"b96b005f",
		16#16ca# => X"bc0b0000",
		16#16cb# => X"1000001d",
		16#16cc# => X"9c21fffc",
		16#16cd# => X"bc05002c",
		16#16ce# => X"100000ba",
		16#16cf# => X"9d600000",
		16#16d0# => X"9de40018",
		16#16d1# => X"9da4000c",
		16#16d2# => X"9d840014",
		16#16d3# => X"9e240010",
		16#16d4# => X"9d040008",
		16#16d5# => X"9e640004",
		16#16d6# => X"18400001",
		16#16d7# => X"b8eb0002",
		16#16d8# => X"a84283b0",
		16#16d9# => X"e0e71000",
		16#16da# => X"84e70000",
		16#16db# => X"44003800",
		16#16dc# => X"15000000",
		16#16dd# => X"9ca5ffd0",
		16#16de# => X"a4a500ff",
		16#16df# => X"bca50009",
		16#16e0# => X"10000015",
		16#16e1# => X"9ca00001",
		16#16e2# => X"9c840004",
		16#16e3# => X"84a40000",
		16#16e4# => X"9ca50001",
		16#16e5# => X"d4042800",
		16#16e6# => X"9cc60001",
		16#16e7# => X"9d600001",
		16#16e8# => X"9c210004",
		16#16e9# => X"d4033000",
		16#16ea# => X"44004800",
		16#16eb# => X"8441fffc",
		16#16ec# => X"9ca5ffd0",
		16#16ed# => X"a4a500ff",
		16#16ee# => X"bc450009",
		16#16ef# => X"10000070",
		16#16f0# => X"9ca00001",
		16#16f1# => X"84ef0000",
		16#16f2# => X"9d600007",
		16#16f3# => X"e0e72800",
		16#16f4# => X"d40f3800",
		16#16f5# => X"9cc60001",
		16#16f6# => X"bc050000",
		16#16f7# => X"13fffff1",
		16#16f8# => X"8ca60000",
		16#16f9# => X"bc250000",
		16#16fa# => X"0fffffee",
		16#16fb# => X"bc25002c",
		16#16fc# => X"13ffffda",
		16#16fd# => X"15000000",
		16#16fe# => X"9cc60001",
		16#16ff# => X"9c210004",
		16#1700# => X"d4033000",
		16#1701# => X"44004800",
		16#1702# => X"8441fffc",
		16#1703# => X"ace50065",
		16#1704# => X"9ce7ffff",
		16#1705# => X"bd870000",
		16#1706# => X"1000004d",
		16#1707# => X"ace50045",
		16#1708# => X"9ce7ffff",
		16#1709# => X"bd670000",
		16#170a# => X"0c000049",
		16#170b# => X"15000000",
		16#170c# => X"9ca5ffd0",
		16#170d# => X"a4a500ff",
		16#170e# => X"bca50009",
		16#170f# => X"13ffffe6",
		16#1710# => X"9ca00001",
		16#1711# => X"9c840014",
		16#1712# => X"84a40000",
		16#1713# => X"9ca50001",
		16#1714# => X"03ffffd2",
		16#1715# => X"d4042800",
		16#1716# => X"9ce5ffd0",
		16#1717# => X"a4e700ff",
		16#1718# => X"bc470009",
		16#1719# => X"1000004b",
		16#171a# => X"bc25002e",
		16#171b# => X"84e80000",
		16#171c# => X"9ca00001",
		16#171d# => X"9d600004",
		16#171e# => X"e0e72800",
		16#171f# => X"03ffffd6",
		16#1720# => X"d4083800",
		16#1721# => X"bc25002e",
		16#1722# => X"0c00005b",
		16#1723# => X"15000000",
		16#1724# => X"9ca5ffd0",
		16#1725# => X"a4a500ff",
		16#1726# => X"bca50009",
		16#1727# => X"13ffffce",
		16#1728# => X"9ca00001",
		16#1729# => X"9c840010",
		16#172a# => X"84a40000",
		16#172b# => X"9ca50001",
		16#172c# => X"03ffffba",
		16#172d# => X"d4042800",
		16#172e# => X"acab0001",
		16#172f# => X"e0a02802",
		16#1730# => X"03ffffc5",
		16#1731# => X"b8a5005f",
		16#1732# => X"9ce5ffd0",
		16#1733# => X"a4e700ff",
		16#1734# => X"bca70009",
		16#1735# => X"10000008",
		16#1736# => X"9d600004",
		16#1737# => X"ace5002d",
		16#1738# => X"9ce7ffff",
		16#1739# => X"bd870000",
		16#173a# => X"0c000031",
		16#173b# => X"ace5002b",
		16#173c# => X"9d600002",
		16#173d# => X"84e40000",
		16#173e# => X"acab0001",
		16#173f# => X"9ce70001",
		16#1740# => X"e0a02802",
		16#1741# => X"d4043800",
		16#1742# => X"03ffffb3",
		16#1743# => X"b8a5005f",
		16#1744# => X"ace5002d",
		16#1745# => X"9ce7ffff",
		16#1746# => X"bd870000",
		16#1747# => X"10000012",
		16#1748# => X"15000000",
		16#1749# => X"aca5002b",
		16#174a# => X"9ca5ffff",
		16#174b# => X"bd650000",
		16#174c# => X"0c00000d",
		16#174d# => X"15000000",
		16#174e# => X"9c84000c",
		16#174f# => X"84a40000",
		16#1750# => X"9ca50001",
		16#1751# => X"03ffff95",
		16#1752# => X"d4042800",
		16#1753# => X"84ec0000",
		16#1754# => X"9ca00001",
		16#1755# => X"9d600003",
		16#1756# => X"e0e72800",
		16#1757# => X"03ffff9e",
		16#1758# => X"d40c3800",
		16#1759# => X"84ed0000",
		16#175a# => X"9ca00001",
		16#175b# => X"9d600006",
		16#175c# => X"e0e72800",
		16#175d# => X"03ffff98",
		16#175e# => X"d40d3800",
		16#175f# => X"9c840018",
		16#1760# => X"84a40000",
		16#1761# => X"9ca50001",
		16#1762# => X"03ffff84",
		16#1763# => X"d4042800",
		16#1764# => X"0c00001f",
		16#1765# => X"9ca00001",
		16#1766# => X"9c840008",
		16#1767# => X"84a40000",
		16#1768# => X"9ca50001",
		16#1769# => X"03ffff7d",
		16#176a# => X"d4042800",
		16#176b# => X"9ce7ffff",
		16#176c# => X"bd870000",
		16#176d# => X"13ffffd0",
		16#176e# => X"9d600002",
		16#176f# => X"bc05002e",
		16#1770# => X"13ffffcd",
		16#1771# => X"9d600005",
		16#1772# => X"84b30000",
		16#1773# => X"9d600001",
		16#1774# => X"e0a55800",
		16#1775# => X"d4132800",
		16#1776# => X"acab0001",
		16#1777# => X"84e40000",
		16#1778# => X"e0a02802",
		16#1779# => X"9ce70001",
		16#177a# => X"b8a5005f",
		16#177b# => X"03ffff7a",
		16#177c# => X"d4043800",
		16#177d# => X"84f10000",
		16#177e# => X"9ca00001",
		16#177f# => X"9d600005",
		16#1780# => X"e0e72800",
		16#1781# => X"03ffff74",
		16#1782# => X"d4113800",
		16#1783# => X"84e80000",
		16#1784# => X"9d600005",
		16#1785# => X"e0e72800",
		16#1786# => X"03ffff6f",
		16#1787# => X"d4083800",
		16#1788# => X"03ffff77",
		16#1789# => X"9cc60001",
		16#178a# => X"d7e117dc",
		16#178b# => X"d7e177e0",
		16#178c# => X"d7e1a7ec",
		16#178d# => X"d7e1b7f0",
		16#178e# => X"d7e1c7f4",
		16#178f# => X"d7e1d7f8",
		16#1790# => X"a8440000",
		16#1791# => X"d7e14ffc",
		16#1792# => X"9c800000",
		16#1793# => X"d7e187e4",
		16#1794# => X"d7e197e8",
		16#1795# => X"9c21ff98",
		16#1796# => X"b8a50010",
		16#1797# => X"d4012000",
		16#1798# => X"d4011040",
		16#1799# => X"d4012020",
		16#179a# => X"d4012004",
		16#179b# => X"d4012024",
		16#179c# => X"d4012008",
		16#179d# => X"d4012028",
		16#179e# => X"d401200c",
		16#179f# => X"d401202c",
		16#17a0# => X"d4012010",
		16#17a1# => X"d4012030",
		16#17a2# => X"d4012014",
		16#17a3# => X"d4012034",
		16#17a4# => X"d4012018",
		16#17a5# => X"d4012038",
		16#17a6# => X"d401201c",
		16#17a7# => X"d401203c",
		16#17a8# => X"b8c60010",
		16#17a9# => X"8d620000",
		16#17aa# => X"b8e70010",
		16#17ab# => X"a9c30000",
		16#17ac# => X"bb050090",
		16#17ad# => X"bac60090",
		16#17ae# => X"ba870090",
		16#17af# => X"e40b2000",
		16#17b0# => X"10000013",
		16#17b1# => X"a748ffff",
		16#17b2# => X"9e410040",
		16#17b3# => X"a8720000",
		16#17b4# => X"07ffff11",
		16#17b5# => X"a8810000",
		16#17b6# => X"b96b0002",
		16#17b7# => X"9c610044",
		16#17b8# => X"e0a35800",
		16#17b9# => X"9ca5ffdc",
		16#17ba# => X"84c50000",
		16#17bb# => X"9cc60001",
		16#17bc# => X"d4053000",
		16#17bd# => X"84a10040",
		16#17be# => X"8ca50000",
		16#17bf# => X"bc250000",
		16#17c0# => X"13fffff4",
		16#17c1# => X"a8720000",
		16#17c2# => X"8d620000",
		16#17c3# => X"e1c27000",
		16#17c4# => X"e4627000",
		16#17c5# => X"10000011",
		16#17c6# => X"d4011040",
		16#17c7# => X"a8a20000",
		16#17c8# => X"00000004",
		16#17c9# => X"a8c20000",
		16#17ca# => X"8d650000",
		16#17cb# => X"a8c50000",
		16#17cc# => X"bc0b002c",
		16#17cd# => X"10000004",
		16#17ce# => X"e06bc005",
		16#17cf# => X"d8061800",
		16#17d0# => X"84a10040",
		16#17d1# => X"e0a5a000",
		16#17d2# => X"e4657000",
		16#17d3# => X"0ffffff7",
		16#17d4# => X"d4012840",
		16#17d5# => X"8d620000",
		16#17d6# => X"bc0b0000",
		16#17d7# => X"10000012",
		16#17d8# => X"d4011040",
		16#17d9# => X"9e410040",
		16#17da# => X"a8720000",
		16#17db# => X"07fffeea",
		16#17dc# => X"a8810000",
		16#17dd# => X"b96b0002",
		16#17de# => X"9c810044",
		16#17df# => X"e0a45800",
		16#17e0# => X"9ca5ffdc",
		16#17e1# => X"84650000",
		16#17e2# => X"9c630001",
		16#17e3# => X"d4051800",
		16#17e4# => X"84610040",
		16#17e5# => X"8c630000",
		16#17e6# => X"bc230000",
		16#17e7# => X"13fffff4",
		16#17e8# => X"a8720000",
		16#17e9# => X"e4627000",
		16#17ea# => X"1000000e",
		16#17eb# => X"d4011040",
		16#17ec# => X"a8a20000",
		16#17ed# => X"8c620000",
		16#17ee# => X"bc03002c",
		16#17ef# => X"10000004",
		16#17f0# => X"e0c3b005",
		16#17f1# => X"d8023000",
		16#17f2# => X"84a10040",
		16#17f3# => X"e045a000",
		16#17f4# => X"d4011040",
		16#17f5# => X"e4827000",
		16#17f6# => X"13fffff7",
		16#17f7# => X"a8a20000",
		16#17f8# => X"84610020",
		16#17f9# => X"04000176",
		16#17fa# => X"a89a0000",
		16#17fb# => X"84610000",
		16#17fc# => X"04000173",
		16#17fd# => X"a88b0000",
		16#17fe# => X"84610024",
		16#17ff# => X"04000170",
		16#1800# => X"a88b0000",
		16#1801# => X"84610004",
		16#1802# => X"0400016d",
		16#1803# => X"a88b0000",
		16#1804# => X"84610028",
		16#1805# => X"0400016a",
		16#1806# => X"a88b0000",
		16#1807# => X"84610008",
		16#1808# => X"04000167",
		16#1809# => X"a88b0000",
		16#180a# => X"8461002c",
		16#180b# => X"04000164",
		16#180c# => X"a88b0000",
		16#180d# => X"8461000c",
		16#180e# => X"04000161",
		16#180f# => X"a88b0000",
		16#1810# => X"84610030",
		16#1811# => X"0400015e",
		16#1812# => X"a88b0000",
		16#1813# => X"84610010",
		16#1814# => X"0400015b",
		16#1815# => X"a88b0000",
		16#1816# => X"84610034",
		16#1817# => X"04000158",
		16#1818# => X"a88b0000",
		16#1819# => X"84610014",
		16#181a# => X"04000155",
		16#181b# => X"a88b0000",
		16#181c# => X"84610038",
		16#181d# => X"04000152",
		16#181e# => X"a88b0000",
		16#181f# => X"84610018",
		16#1820# => X"0400014f",
		16#1821# => X"a88b0000",
		16#1822# => X"8461003c",
		16#1823# => X"0400014c",
		16#1824# => X"a88b0000",
		16#1825# => X"8461001c",
		16#1826# => X"04000149",
		16#1827# => X"a88b0000",
		16#1828# => X"9c210068",
		16#1829# => X"8521fffc",
		16#182a# => X"8441ffdc",
		16#182b# => X"85c1ffe0",
		16#182c# => X"8601ffe4",
		16#182d# => X"8641ffe8",
		16#182e# => X"8681ffec",
		16#182f# => X"86c1fff0",
		16#1830# => X"8701fff4",
		16#1831# => X"44004800",
		16#1832# => X"8741fff8",
		16#1833# => X"d7e117fc",
		16#1834# => X"bc430005",
		16#1835# => X"0c000006",
		16#1836# => X"9c21fffc",
		16#1837# => X"9c210004",
		16#1838# => X"9d600000",
		16#1839# => X"44004800",
		16#183a# => X"8441fffc",
		16#183b# => X"18400001",
		16#183c# => X"b8630002",
		16#183d# => X"a8428490",
		16#183e# => X"e0631000",
		16#183f# => X"84630000",
		16#1840# => X"44001800",
		16#1841# => X"15000000",
		16#1842# => X"18600001",
		16#1843# => X"a863b800",
		16#1844# => X"85630000",
		16#1845# => X"9c210004",
		16#1846# => X"44004800",
		16#1847# => X"8441fffc",
		16#1848# => X"18600001",
		16#1849# => X"a863b804",
		16#184a# => X"85630000",
		16#184b# => X"9c210004",
		16#184c# => X"44004800",
		16#184d# => X"8441fffc",
		16#184e# => X"18600001",
		16#184f# => X"a863add8",
		16#1850# => X"85630000",
		16#1851# => X"9c210004",
		16#1852# => X"44004800",
		16#1853# => X"8441fffc",
		16#1854# => X"18600001",
		16#1855# => X"a863addc",
		16#1856# => X"85630000",
		16#1857# => X"9c210004",
		16#1858# => X"44004800",
		16#1859# => X"8441fffc",
		16#185a# => X"18600001",
		16#185b# => X"a863b808",
		16#185c# => X"85630000",
		16#185d# => X"9c210004",
		16#185e# => X"44004800",
		16#185f# => X"8441fffc",
		16#1860# => X"a484ffff",
		16#1861# => X"a46300ff",
		16#1862# => X"ace44002",
		16#1863# => X"e0c32005",
		16#1864# => X"b8e70041",
		16#1865# => X"a4c60001",
		16#1866# => X"b8a30041",
		16#1867# => X"a8e78000",
		16#1868# => X"bc260001",
		16#1869# => X"0c000041",
		16#186a# => X"b8640041",
		16#186b# => X"ace34002",
		16#186c# => X"e0c51805",
		16#186d# => X"b8e70041",
		16#186e# => X"a4c60001",
		16#186f# => X"b8850041",
		16#1870# => X"a8e78000",
		16#1871# => X"bc260001",
		16#1872# => X"0c000047",
		16#1873# => X"b8630041",
		16#1874# => X"acc34002",
		16#1875# => X"e0a41805",
		16#1876# => X"b8c60041",
		16#1877# => X"a4a50001",
		16#1878# => X"b8840041",
		16#1879# => X"a8c68000",
		16#187a# => X"bc250001",
		16#187b# => X"0c00003c",
		16#187c# => X"b8630041",
		16#187d# => X"acc34002",
		16#187e# => X"e0a41805",
		16#187f# => X"b8c60041",
		16#1880# => X"a4a50001",
		16#1881# => X"b8840041",
		16#1882# => X"a8c68000",
		16#1883# => X"bc250001",
		16#1884# => X"0c000031",
		16#1885# => X"b8630041",
		16#1886# => X"acc34002",
		16#1887# => X"e0a41805",
		16#1888# => X"b8c60041",
		16#1889# => X"a4a50001",
		16#188a# => X"b8840041",
		16#188b# => X"a8c68000",
		16#188c# => X"bc250001",
		16#188d# => X"0c000026",
		16#188e# => X"b8630041",
		16#188f# => X"acc34002",
		16#1890# => X"e0a41805",
		16#1891# => X"b8c60041",
		16#1892# => X"a4a50001",
		16#1893# => X"b8840041",
		16#1894# => X"a8c68000",
		16#1895# => X"bc250001",
		16#1896# => X"0c00001b",
		16#1897# => X"b8630041",
		16#1898# => X"acc34002",
		16#1899# => X"e0a41805",
		16#189a# => X"b8c60041",
		16#189b# => X"a4a50001",
		16#189c# => X"b8630041",
		16#189d# => X"bc250001",
		16#189e# => X"0c000011",
		16#189f# => X"a8c68000",
		16#18a0# => X"acc34002",
		16#18a1# => X"b8840041",
		16#18a2# => X"b8c60041",
		16#18a3# => X"a4a30001",
		16#18a4# => X"b8630041",
		16#18a5# => X"e4052000",
		16#18a6# => X"0c000006",
		16#18a7# => X"a8c68000",
		16#18a8# => X"44004800",
		16#18a9# => X"a563ffff",
		16#18aa# => X"03ffffc1",
		16#18ab# => X"a8670000",
		16#18ac# => X"a8660000",
		16#18ad# => X"44004800",
		16#18ae# => X"a563ffff",
		16#18af# => X"03fffff1",
		16#18b0# => X"a8660000",
		16#18b1# => X"03ffffe7",
		16#18b2# => X"a8660000",
		16#18b3# => X"03ffffdc",
		16#18b4# => X"a8660000",
		16#18b5# => X"03ffffd1",
		16#18b6# => X"a8660000",
		16#18b7# => X"03ffffc6",
		16#18b8# => X"a8660000",
		16#18b9# => X"03ffffbb",
		16#18ba# => X"a8670000",
		16#18bb# => X"a463ffff",
		16#18bc# => X"a484ffff",
		16#18bd# => X"a4a300ff",
		16#18be# => X"ace44002",
		16#18bf# => X"e0c52005",
		16#18c0# => X"b8e70041",
		16#18c1# => X"a4c60001",
		16#18c2# => X"b8a50041",
		16#18c3# => X"a8e78000",
		16#18c4# => X"bc260001",
		16#18c5# => X"0c000089",
		16#18c6# => X"b8840041",
		16#18c7# => X"ace44002",
		16#18c8# => X"e0c52005",
		16#18c9# => X"b8e70041",
		16#18ca# => X"a4c60001",
		16#18cb# => X"b8a50041",
		16#18cc# => X"a8e78000",
		16#18cd# => X"bc260001",
		16#18ce# => X"0c00009f",
		16#18cf# => X"b8840041",
		16#18d0# => X"ace44002",
		16#18d1# => X"e0c52005",
		16#18d2# => X"b8e70041",
		16#18d3# => X"a4c60001",
		16#18d4# => X"b8a50041",
		16#18d5# => X"a8e78000",
		16#18d6# => X"bc260001",
		16#18d7# => X"0c000094",
		16#18d8# => X"b8840041",
		16#18d9# => X"ace44002",
		16#18da# => X"e0c52005",
		16#18db# => X"b8e70041",
		16#18dc# => X"a4c60001",
		16#18dd# => X"b8a50041",
		16#18de# => X"a8e78000",
		16#18df# => X"bc260001",
		16#18e0# => X"0c000089",
		16#18e1# => X"b8840041",
		16#18e2# => X"ace44002",
		16#18e3# => X"e0c52005",
		16#18e4# => X"b8e70041",
		16#18e5# => X"a4c60001",
		16#18e6# => X"b8a50041",
		16#18e7# => X"a8e78000",
		16#18e8# => X"bc260001",
		16#18e9# => X"0c00007e",
		16#18ea# => X"b8840041",
		16#18eb# => X"ace44002",
		16#18ec# => X"e0c52005",
		16#18ed# => X"b8e70041",
		16#18ee# => X"a4c60001",
		16#18ef# => X"b8a50041",
		16#18f0# => X"a8e78000",
		16#18f1# => X"bc260001",
		16#18f2# => X"0c000073",
		16#18f3# => X"b8840041",
		16#18f4# => X"ace44002",
		16#18f5# => X"e0c52005",
		16#18f6# => X"b8e70041",
		16#18f7# => X"a4c60001",
		16#18f8# => X"b8840041",
		16#18f9# => X"bc260001",
		16#18fa# => X"0c000069",
		16#18fb# => X"a8e78000",
		16#18fc# => X"ace44002",
		16#18fd# => X"b8a50041",
		16#18fe# => X"b8e70041",
		16#18ff# => X"a4c40001",
		16#1900# => X"b8840041",
		16#1901# => X"e4062800",
		16#1902# => X"0c00005f",
		16#1903# => X"a8e78000",
		16#1904# => X"b8a30048",
		16#1905# => X"ace44002",
		16#1906# => X"b8640041",
		16#1907# => X"e0842805",
		16#1908# => X"b8e70041",
		16#1909# => X"a4c40001",
		16#190a# => X"a4a500ff",
		16#190b# => X"a8e78000",
		16#190c# => X"bc260001",
		16#190d# => X"0c000052",
		16#190e# => X"b8850041",
		16#190f# => X"acc34002",
		16#1910# => X"e0a41805",
		16#1911# => X"b8c60041",
		16#1912# => X"a4a50001",
		16#1913# => X"b8840041",
		16#1914# => X"a8c68000",
		16#1915# => X"bc250001",
		16#1916# => X"0c000047",
		16#1917# => X"b8630041",
		16#1918# => X"acc34002",
		16#1919# => X"e0a41805",
		16#191a# => X"b8c60041",
		16#191b# => X"a4a50001",
		16#191c# => X"b8840041",
		16#191d# => X"a8c68000",
		16#191e# => X"bc250001",
		16#191f# => X"0c00003c",
		16#1920# => X"b8630041",
		16#1921# => X"acc34002",
		16#1922# => X"e0a41805",
		16#1923# => X"b8c60041",
		16#1924# => X"a4a50001",
		16#1925# => X"b8840041",
		16#1926# => X"a8c68000",
		16#1927# => X"bc250001",
		16#1928# => X"0c000031",
		16#1929# => X"b8630041",
		16#192a# => X"acc34002",
		16#192b# => X"e0a41805",
		16#192c# => X"b8c60041",
		16#192d# => X"a4a50001",
		16#192e# => X"b8840041",
		16#192f# => X"a8c68000",
		16#1930# => X"bc250001",
		16#1931# => X"0c000026",
		16#1932# => X"b8630041",
		16#1933# => X"acc34002",
		16#1934# => X"e0a41805",
		16#1935# => X"b8c60041",
		16#1936# => X"a4a50001",
		16#1937# => X"b8840041",
		16#1938# => X"a8c68000",
		16#1939# => X"bc250001",
		16#193a# => X"0c00001b",
		16#193b# => X"b8630041",
		16#193c# => X"acc34002",
		16#193d# => X"e0a41805",
		16#193e# => X"b8c60041",
		16#193f# => X"a4a50001",
		16#1940# => X"b8630041",
		16#1941# => X"bc250001",
		16#1942# => X"0c000011",
		16#1943# => X"a8c68000",
		16#1944# => X"acc34002",
		16#1945# => X"b8840041",
		16#1946# => X"b8c60041",
		16#1947# => X"a4a30001",
		16#1948# => X"b8630041",
		16#1949# => X"e4052000",
		16#194a# => X"0c000006",
		16#194b# => X"a8c68000",
		16#194c# => X"44004800",
		16#194d# => X"a563ffff",
		16#194e# => X"03ffff79",
		16#194f# => X"a8870000",
		16#1950# => X"a8660000",
		16#1951# => X"44004800",
		16#1952# => X"a563ffff",
		16#1953# => X"03fffff1",
		16#1954# => X"a8660000",
		16#1955# => X"03ffffe7",
		16#1956# => X"a8660000",
		16#1957# => X"03ffffdc",
		16#1958# => X"a8660000",
		16#1959# => X"03ffffd1",
		16#195a# => X"a8660000",
		16#195b# => X"03ffffc6",
		16#195c# => X"a8660000",
		16#195d# => X"03ffffbb",
		16#195e# => X"a8660000",
		16#195f# => X"03ffffb0",
		16#1960# => X"a8670000",
		16#1961# => X"03ffffa3",
		16#1962# => X"a8870000",
		16#1963# => X"03ffff99",
		16#1964# => X"a8870000",
		16#1965# => X"03ffff8f",
		16#1966# => X"a8870000",
		16#1967# => X"03ffff84",
		16#1968# => X"a8870000",
		16#1969# => X"03ffff79",
		16#196a# => X"a8870000",
		16#196b# => X"03ffff6e",
		16#196c# => X"a8870000",
		16#196d# => X"03ffff63",
		16#196e# => X"a8870000",
		16#196f# => X"a4c3ffff",
		16#1970# => X"a484ffff",
		16#1971# => X"a4a600ff",
		16#1972# => X"ad044002",
		16#1973# => X"e0e42805",
		16#1974# => X"b9080041",
		16#1975# => X"a4e70001",
		16#1976# => X"b8a50041",
		16#1977# => X"a9088000",
		16#1978# => X"bc270001",
		16#1979# => X"0c000119",
		16#197a# => X"b8840041",
		16#197b# => X"ad044002",
		16#197c# => X"e0e52005",
		16#197d# => X"b9080041",
		16#197e# => X"a4e70001",
		16#197f# => X"b8a50041",
		16#1980# => X"a9088000",
		16#1981# => X"bc270001",
		16#1982# => X"0c00014f",
		16#1983# => X"b8840041",
		16#1984# => X"ad044002",
		16#1985# => X"e0e52005",
		16#1986# => X"b9080041",
		16#1987# => X"a4e70001",
		16#1988# => X"b8a50041",
		16#1989# => X"a9088000",
		16#198a# => X"bc270001",
		16#198b# => X"0c000144",
		16#198c# => X"b8840041",
		16#198d# => X"ad044002",
		16#198e# => X"e0e52005",
		16#198f# => X"b9080041",
		16#1990# => X"a4e70001",
		16#1991# => X"b8a50041",
		16#1992# => X"a9088000",
		16#1993# => X"bc270001",
		16#1994# => X"0c000139",
		16#1995# => X"b8840041",
		16#1996# => X"ad044002",
		16#1997# => X"e0e52005",
		16#1998# => X"b9080041",
		16#1999# => X"a4e70001",
		16#199a# => X"b8a50041",
		16#199b# => X"a9088000",
		16#199c# => X"bc270001",
		16#199d# => X"0c00012e",
		16#199e# => X"b8840041",
		16#199f# => X"ad044002",
		16#19a0# => X"e0e52005",
		16#19a1# => X"b9080041",
		16#19a2# => X"a4e70001",
		16#19a3# => X"b8a50041",
		16#19a4# => X"a9088000",
		16#19a5# => X"bc270001",
		16#19a6# => X"0c000123",
		16#19a7# => X"b8840041",
		16#19a8# => X"ad044002",
		16#19a9# => X"e0e52005",
		16#19aa# => X"b9080041",
		16#19ab# => X"a4e70001",
		16#19ac# => X"b8840041",
		16#19ad# => X"bc270001",
		16#19ae# => X"0c000119",
		16#19af# => X"a9088000",
		16#19b0# => X"ad044002",
		16#19b1# => X"b8a50041",
		16#19b2# => X"b9080041",
		16#19b3# => X"a4e40001",
		16#19b4# => X"b8840041",
		16#19b5# => X"e4072800",
		16#19b6# => X"0c00010f",
		16#19b7# => X"a9088000",
		16#19b8# => X"b8c60048",
		16#19b9# => X"ad044002",
		16#19ba# => X"b8a40041",
		16#19bb# => X"e0843005",
		16#19bc# => X"b9080041",
		16#19bd# => X"a4e40001",
		16#19be# => X"a4c600ff",
		16#19bf# => X"a9088000",
		16#19c0# => X"bc270001",
		16#19c1# => X"0c000102",
		16#19c2# => X"b8860041",
		16#19c3# => X"ace54002",
		16#19c4# => X"e0c42805",
		16#19c5# => X"b8e70041",
		16#19c6# => X"a4c60001",
		16#19c7# => X"b8840041",
		16#19c8# => X"a8e78000",
		16#19c9# => X"bc260001",
		16#19ca# => X"0c0000f7",
		16#19cb# => X"b8a50041",
		16#19cc# => X"ace54002",
		16#19cd# => X"e0c42805",
		16#19ce# => X"b8e70041",
		16#19cf# => X"a4c60001",
		16#19d0# => X"b8840041",
		16#19d1# => X"a8e78000",
		16#19d2# => X"bc260001",
		16#19d3# => X"0c0000ec",
		16#19d4# => X"b8a50041",
		16#19d5# => X"ace54002",
		16#19d6# => X"e0c42805",
		16#19d7# => X"b8e70041",
		16#19d8# => X"a4c60001",
		16#19d9# => X"b8840041",
		16#19da# => X"a8e78000",
		16#19db# => X"bc260001",
		16#19dc# => X"0c0000e1",
		16#19dd# => X"b8a50041",
		16#19de# => X"ace54002",
		16#19df# => X"e0c42805",
		16#19e0# => X"b8e70041",
		16#19e1# => X"a4c60001",
		16#19e2# => X"b8840041",
		16#19e3# => X"a8e78000",
		16#19e4# => X"bc260001",
		16#19e5# => X"0c0000d6",
		16#19e6# => X"b8a50041",
		16#19e7# => X"ace54002",
		16#19e8# => X"e0c42805",
		16#19e9# => X"b8e70041",
		16#19ea# => X"a4c60001",
		16#19eb# => X"b8840041",
		16#19ec# => X"a8e78000",
		16#19ed# => X"bc260001",
		16#19ee# => X"0c0000cb",
		16#19ef# => X"b8a50041",
		16#19f0# => X"ace54002",
		16#19f1# => X"e0c42805",
		16#19f2# => X"b8e70041",
		16#19f3# => X"a4c60001",
		16#19f4# => X"b8a50041",
		16#19f5# => X"bc260001",
		16#19f6# => X"0c0000c1",
		16#19f7# => X"a8e78000",
		16#19f8# => X"ace54002",
		16#19f9# => X"b8840041",
		16#19fa# => X"b8e70041",
		16#19fb# => X"a4c50001",
		16#19fc# => X"b8a50041",
		16#19fd# => X"e4062000",
		16#19fe# => X"0c0000b7",
		16#19ff# => X"a8e78000",
		16#1a00# => X"b8630050",
		16#1a01# => X"ace54002",
		16#1a02# => X"b8850041",
		16#1a03# => X"a4c300ff",
		16#1a04# => X"b8e70041",
		16#1a05# => X"e1062805",
		16#1a06# => X"b8a60041",
		16#1a07# => X"a4c80001",
		16#1a08# => X"bc260001",
		16#1a09# => X"0c0000aa",
		16#1a0a# => X"a8e78000",
		16#1a0b# => X"ace44002",
		16#1a0c# => X"e0c52005",
		16#1a0d# => X"b8e70041",
		16#1a0e# => X"a4c60001",
		16#1a0f# => X"b8a50041",
		16#1a10# => X"a8e78000",
		16#1a11# => X"bc260001",
		16#1a12# => X"0c00009f",
		16#1a13# => X"b8840041",
		16#1a14# => X"ace44002",
		16#1a15# => X"e0c52005",
		16#1a16# => X"b8e70041",
		16#1a17# => X"a4c60001",
		16#1a18# => X"b8a50041",
		16#1a19# => X"a8e78000",
		16#1a1a# => X"bc260001",
		16#1a1b# => X"0c000094",
		16#1a1c# => X"b8840041",
		16#1a1d# => X"ace44002",
		16#1a1e# => X"e0c52005",
		16#1a1f# => X"b8e70041",
		16#1a20# => X"a4c60001",
		16#1a21# => X"b8a50041",
		16#1a22# => X"a8e78000",
		16#1a23# => X"bc260001",
		16#1a24# => X"0c000089",
		16#1a25# => X"b8840041",
		16#1a26# => X"ace44002",
		16#1a27# => X"e0c52005",
		16#1a28# => X"b8e70041",
		16#1a29# => X"a4c60001",
		16#1a2a# => X"b8a50041",
		16#1a2b# => X"a8e78000",
		16#1a2c# => X"bc260001",
		16#1a2d# => X"0c00007e",
		16#1a2e# => X"b8840041",
		16#1a2f# => X"ace44002",
		16#1a30# => X"e0c52005",
		16#1a31# => X"b8e70041",
		16#1a32# => X"a4c60001",
		16#1a33# => X"b8a50041",
		16#1a34# => X"a8e78000",
		16#1a35# => X"bc260001",
		16#1a36# => X"0c000073",
		16#1a37# => X"b8840041",
		16#1a38# => X"ace44002",
		16#1a39# => X"e0c52005",
		16#1a3a# => X"b8e70041",
		16#1a3b# => X"a4c60001",
		16#1a3c# => X"b8840041",
		16#1a3d# => X"bc260001",
		16#1a3e# => X"0c000069",
		16#1a3f# => X"a8e78000",
		16#1a40# => X"ace44002",
		16#1a41# => X"b8a50041",
		16#1a42# => X"b8e70041",
		16#1a43# => X"a4c40001",
		16#1a44# => X"b8840041",
		16#1a45# => X"e4062800",
		16#1a46# => X"0c00005f",
		16#1a47# => X"a8e78000",
		16#1a48# => X"b8a30048",
		16#1a49# => X"ace44002",
		16#1a4a# => X"b8640041",
		16#1a4b# => X"e0842805",
		16#1a4c# => X"b8e70041",
		16#1a4d# => X"a4c40001",
		16#1a4e# => X"a4a500ff",
		16#1a4f# => X"a8e78000",
		16#1a50# => X"bc260001",
		16#1a51# => X"0c000052",
		16#1a52# => X"b8850041",
		16#1a53# => X"acc34002",
		16#1a54# => X"e0a41805",
		16#1a55# => X"b8c60041",
		16#1a56# => X"a4a50001",
		16#1a57# => X"b8840041",
		16#1a58# => X"a8c68000",
		16#1a59# => X"bc250001",
		16#1a5a# => X"0c000047",
		16#1a5b# => X"b8630041",
		16#1a5c# => X"acc34002",
		16#1a5d# => X"e0a41805",
		16#1a5e# => X"b8c60041",
		16#1a5f# => X"a4a50001",
		16#1a60# => X"b8840041",
		16#1a61# => X"a8c68000",
		16#1a62# => X"bc250001",
		16#1a63# => X"0c00003c",
		16#1a64# => X"b8630041",
		16#1a65# => X"acc34002",
		16#1a66# => X"e0a41805",
		16#1a67# => X"b8c60041",
		16#1a68# => X"a4a50001",
		16#1a69# => X"b8840041",
		16#1a6a# => X"a8c68000",
		16#1a6b# => X"bc250001",
		16#1a6c# => X"0c000031",
		16#1a6d# => X"b8630041",
		16#1a6e# => X"acc34002",
		16#1a6f# => X"e0a41805",
		16#1a70# => X"b8c60041",
		16#1a71# => X"a4a50001",
		16#1a72# => X"b8840041",
		16#1a73# => X"a8c68000",
		16#1a74# => X"bc250001",
		16#1a75# => X"0c000026",
		16#1a76# => X"b8630041",
		16#1a77# => X"acc34002",
		16#1a78# => X"e0a41805",
		16#1a79# => X"b8c60041",
		16#1a7a# => X"a4a50001",
		16#1a7b# => X"b8840041",
		16#1a7c# => X"a8c68000",
		16#1a7d# => X"bc250001",
		16#1a7e# => X"0c00001b",
		16#1a7f# => X"b8630041",
		16#1a80# => X"acc34002",
		16#1a81# => X"e0a41805",
		16#1a82# => X"b8c60041",
		16#1a83# => X"a4a50001",
		16#1a84# => X"b8630041",
		16#1a85# => X"bc250001",
		16#1a86# => X"0c000011",
		16#1a87# => X"a8c68000",
		16#1a88# => X"acc34002",
		16#1a89# => X"b8840041",
		16#1a8a# => X"b8c60041",
		16#1a8b# => X"a4a30001",
		16#1a8c# => X"b8630041",
		16#1a8d# => X"e4052000",
		16#1a8e# => X"0c000006",
		16#1a8f# => X"a8c68000",
		16#1a90# => X"44004800",
		16#1a91# => X"a563ffff",
		16#1a92# => X"03fffee9",
		16#1a93# => X"a8880000",
		16#1a94# => X"a8660000",
		16#1a95# => X"44004800",
		16#1a96# => X"a563ffff",
		16#1a97# => X"03fffff1",
		16#1a98# => X"a8660000",
		16#1a99# => X"03ffffe7",
		16#1a9a# => X"a8660000",
		16#1a9b# => X"03ffffdc",
		16#1a9c# => X"a8660000",
		16#1a9d# => X"03ffffd1",
		16#1a9e# => X"a8660000",
		16#1a9f# => X"03ffffc6",
		16#1aa0# => X"a8660000",
		16#1aa1# => X"03ffffbb",
		16#1aa2# => X"a8660000",
		16#1aa3# => X"03ffffb0",
		16#1aa4# => X"a8670000",
		16#1aa5# => X"03ffffa3",
		16#1aa6# => X"a8870000",
		16#1aa7# => X"03ffff99",
		16#1aa8# => X"a8870000",
		16#1aa9# => X"03ffff8f",
		16#1aaa# => X"a8870000",
		16#1aab# => X"03ffff84",
		16#1aac# => X"a8870000",
		16#1aad# => X"03ffff79",
		16#1aae# => X"a8870000",
		16#1aaf# => X"03ffff6e",
		16#1ab0# => X"a8870000",
		16#1ab1# => X"03ffff63",
		16#1ab2# => X"a8870000",
		16#1ab3# => X"03ffff58",
		16#1ab4# => X"a8870000",
		16#1ab5# => X"03ffff4b",
		16#1ab6# => X"a8a70000",
		16#1ab7# => X"03ffff41",
		16#1ab8# => X"a8a70000",
		16#1ab9# => X"03ffff37",
		16#1aba# => X"a8a70000",
		16#1abb# => X"03ffff2c",
		16#1abc# => X"a8a70000",
		16#1abd# => X"03ffff21",
		16#1abe# => X"a8a70000",
		16#1abf# => X"03ffff16",
		16#1ac0# => X"a8a70000",
		16#1ac1# => X"03ffff0b",
		16#1ac2# => X"a8a70000",
		16#1ac3# => X"03ffff00",
		16#1ac4# => X"a8a80000",
		16#1ac5# => X"03fffef3",
		16#1ac6# => X"a8880000",
		16#1ac7# => X"03fffee9",
		16#1ac8# => X"a8880000",
		16#1ac9# => X"03fffedf",
		16#1aca# => X"a8880000",
		16#1acb# => X"03fffed4",
		16#1acc# => X"a8880000",
		16#1acd# => X"03fffec9",
		16#1ace# => X"a8880000",
		16#1acf# => X"03fffebe",
		16#1ad0# => X"a8880000",
		16#1ad1# => X"03fffeb3",
		16#1ad2# => X"a8880000",
		16#1ad3# => X"a463ffff",
		16#1ad4# => X"a484ffff",
		16#1ad5# => X"a4a300ff",
		16#1ad6# => X"ace44002",
		16#1ad7# => X"e0c42805",
		16#1ad8# => X"b8e70041",
		16#1ad9# => X"a4c60001",
		16#1ada# => X"b8a50041",
		16#1adb# => X"a8e78000",
		16#1adc# => X"bc260001",
		16#1add# => X"0c000089",
		16#1ade# => X"b8840041",
		16#1adf# => X"ace44002",
		16#1ae0# => X"e0c52005",
		16#1ae1# => X"b8e70041",
		16#1ae2# => X"a4c60001",
		16#1ae3# => X"b8a50041",
		16#1ae4# => X"a8e78000",
		16#1ae5# => X"bc260001",
		16#1ae6# => X"0c00009f",
		16#1ae7# => X"b8840041",
		16#1ae8# => X"ace44002",
		16#1ae9# => X"e0c52005",
		16#1aea# => X"b8e70041",
		16#1aeb# => X"a4c60001",
		16#1aec# => X"b8a50041",
		16#1aed# => X"a8e78000",
		16#1aee# => X"bc260001",
		16#1aef# => X"0c000094",
		16#1af0# => X"b8840041",
		16#1af1# => X"ace44002",
		16#1af2# => X"e0c52005",
		16#1af3# => X"b8e70041",
		16#1af4# => X"a4c60001",
		16#1af5# => X"b8a50041",
		16#1af6# => X"a8e78000",
		16#1af7# => X"bc260001",
		16#1af8# => X"0c000089",
		16#1af9# => X"b8840041",
		16#1afa# => X"ace44002",
		16#1afb# => X"e0c52005",
		16#1afc# => X"b8e70041",
		16#1afd# => X"a4c60001",
		16#1afe# => X"b8a50041",
		16#1aff# => X"a8e78000",
		16#1b00# => X"bc260001",
		16#1b01# => X"0c00007e",
		16#1b02# => X"b8840041",
		16#1b03# => X"ace44002",
		16#1b04# => X"e0c52005",
		16#1b05# => X"b8e70041",
		16#1b06# => X"a4c60001",
		16#1b07# => X"b8a50041",
		16#1b08# => X"a8e78000",
		16#1b09# => X"bc260001",
		16#1b0a# => X"0c000073",
		16#1b0b# => X"b8840041",
		16#1b0c# => X"ace44002",
		16#1b0d# => X"e0c52005",
		16#1b0e# => X"b8e70041",
		16#1b0f# => X"a4c60001",
		16#1b10# => X"b8840041",
		16#1b11# => X"bc260001",
		16#1b12# => X"0c000069",
		16#1b13# => X"a8e78000",
		16#1b14# => X"ace44002",
		16#1b15# => X"b8a50041",
		16#1b16# => X"b8e70041",
		16#1b17# => X"a4c40001",
		16#1b18# => X"b8840041",
		16#1b19# => X"e4062800",
		16#1b1a# => X"0c00005f",
		16#1b1b# => X"a8e78000",
		16#1b1c# => X"b8a30048",
		16#1b1d# => X"ace44002",
		16#1b1e# => X"b8640041",
		16#1b1f# => X"e0842805",
		16#1b20# => X"b8e70041",
		16#1b21# => X"a4c40001",
		16#1b22# => X"a4a500ff",
		16#1b23# => X"a8e78000",
		16#1b24# => X"bc260001",
		16#1b25# => X"0c000052",
		16#1b26# => X"b8850041",
		16#1b27# => X"acc34002",
		16#1b28# => X"e0a41805",
		16#1b29# => X"b8c60041",
		16#1b2a# => X"a4a50001",
		16#1b2b# => X"b8840041",
		16#1b2c# => X"a8c68000",
		16#1b2d# => X"bc250001",
		16#1b2e# => X"0c000047",
		16#1b2f# => X"b8630041",
		16#1b30# => X"acc34002",
		16#1b31# => X"e0a41805",
		16#1b32# => X"b8c60041",
		16#1b33# => X"a4a50001",
		16#1b34# => X"b8840041",
		16#1b35# => X"a8c68000",
		16#1b36# => X"bc250001",
		16#1b37# => X"0c00003c",
		16#1b38# => X"b8630041",
		16#1b39# => X"acc34002",
		16#1b3a# => X"e0a41805",
		16#1b3b# => X"b8c60041",
		16#1b3c# => X"a4a50001",
		16#1b3d# => X"b8840041",
		16#1b3e# => X"a8c68000",
		16#1b3f# => X"bc250001",
		16#1b40# => X"0c000031",
		16#1b41# => X"b8630041",
		16#1b42# => X"acc34002",
		16#1b43# => X"e0a41805",
		16#1b44# => X"b8c60041",
		16#1b45# => X"a4a50001",
		16#1b46# => X"b8840041",
		16#1b47# => X"a8c68000",
		16#1b48# => X"bc250001",
		16#1b49# => X"0c000026",
		16#1b4a# => X"b8630041",
		16#1b4b# => X"acc34002",
		16#1b4c# => X"e0a41805",
		16#1b4d# => X"b8c60041",
		16#1b4e# => X"a4a50001",
		16#1b4f# => X"b8840041",
		16#1b50# => X"a8c68000",
		16#1b51# => X"bc250001",
		16#1b52# => X"0c00001b",
		16#1b53# => X"b8630041",
		16#1b54# => X"acc34002",
		16#1b55# => X"e0a41805",
		16#1b56# => X"b8c60041",
		16#1b57# => X"a4a50001",
		16#1b58# => X"b8630041",
		16#1b59# => X"bc250001",
		16#1b5a# => X"0c000011",
		16#1b5b# => X"a8c68000",
		16#1b5c# => X"acc34002",
		16#1b5d# => X"b8840041",
		16#1b5e# => X"b8c60041",
		16#1b5f# => X"a4a30001",
		16#1b60# => X"b8630041",
		16#1b61# => X"e4052000",
		16#1b62# => X"0c000006",
		16#1b63# => X"a8c68000",
		16#1b64# => X"44004800",
		16#1b65# => X"a563ffff",
		16#1b66# => X"03ffff79",
		16#1b67# => X"a8870000",
		16#1b68# => X"a8660000",
		16#1b69# => X"44004800",
		16#1b6a# => X"a563ffff",
		16#1b6b# => X"03fffff1",
		16#1b6c# => X"a8660000",
		16#1b6d# => X"03ffffe7",
		16#1b6e# => X"a8660000",
		16#1b6f# => X"03ffffdc",
		16#1b70# => X"a8660000",
		16#1b71# => X"03ffffd1",
		16#1b72# => X"a8660000",
		16#1b73# => X"03ffffc6",
		16#1b74# => X"a8660000",
		16#1b75# => X"03ffffbb",
		16#1b76# => X"a8660000",
		16#1b77# => X"03ffffb0",
		16#1b78# => X"a8670000",
		16#1b79# => X"03ffffa3",
		16#1b7a# => X"a8870000",
		16#1b7b# => X"03ffff99",
		16#1b7c# => X"a8870000",
		16#1b7d# => X"03ffff8f",
		16#1b7e# => X"a8870000",
		16#1b7f# => X"03ffff84",
		16#1b80# => X"a8870000",
		16#1b81# => X"03ffff79",
		16#1b82# => X"a8870000",
		16#1b83# => X"03ffff6e",
		16#1b84# => X"a8870000",
		16#1b85# => X"03ffff63",
		16#1b86# => X"a8870000",
		16#1b87# => X"44004800",
		16#1b88# => X"9d600000",
		16#1b89# => X"d7e14ffc",
		16#1b8a# => X"040015ec",
		16#1b8b# => X"9c21fff8",
		16#1b8c# => X"bc2b0000",
		16#1b8d# => X"0c000006",
		16#1b8e# => X"15000000",
		16#1b8f# => X"9c210008",
		16#1b90# => X"8521fffc",
		16#1b91# => X"44004800",
		16#1b92# => X"15000000",
		16#1b93# => X"04000a06",
		16#1b94# => X"15000000",
		16#1b95# => X"bc0b0000",
		16#1b96# => X"0c00000d",
		16#1b97# => X"15000000",
		16#1b98# => X"04000a01",
		16#1b99# => X"15000000",
		16#1b9a# => X"18600001",
		16#1b9b# => X"d4015800",
		16#1b9c# => X"040019e2",
		16#1b9d# => X"a8637ebc",
		16#1b9e# => X"18600001",
		16#1b9f# => X"04001ac2",
		16#1ba0# => X"a86384a8",
		16#1ba1# => X"040015c4",
		16#1ba2# => X"9c600001",
		16#1ba3# => X"040009f6",
		16#1ba4# => X"15000000",
		16#1ba5# => X"040009fa",
		16#1ba6# => X"9c6bffff",
		16#1ba7# => X"03fffff1",
		16#1ba8# => X"15000000",
		16#1ba9# => X"d7e14ffc",
		16#1baa# => X"9c21fffc",
		16#1bab# => X"9c210004",
		16#1bac# => X"8521fffc",
		16#1bad# => X"000015d3",
		16#1bae# => X"15000000",
		16#1baf# => X"1860017d",
		16#1bb0# => X"d7e14ffc",
		16#1bb1# => X"a8637840",
		16#1bb2# => X"040000f4",
		16#1bb3# => X"9c21fffc",
		16#1bb4# => X"040009e5",
		16#1bb5# => X"15000000",
		16#1bb6# => X"1860f000",
		16#1bb7# => X"040000f3",
		16#1bb8# => X"a88b0000",
		16#1bb9# => X"040009e0",
		16#1bba# => X"15000000",
		16#1bbb# => X"1860f000",
		16#1bbc# => X"040000f4",
		16#1bbd# => X"a88b0000",
		16#1bbe# => X"040009db",
		16#1bbf# => X"15000000",
		16#1bc0# => X"18a00001",
		16#1bc1# => X"9c210004",
		16#1bc2# => X"1860f000",
		16#1bc3# => X"a88b0000",
		16#1bc4# => X"8521fffc",
		16#1bc5# => X"00000139",
		16#1bc6# => X"a8a5b83c",
		16#1bc7# => X"d7e14ffc",
		16#1bc8# => X"040009d1",
		16#1bc9# => X"9c21fffc",
		16#1bca# => X"18a00001",
		16#1bcb# => X"9c210004",
		16#1bcc# => X"1860f000",
		16#1bcd# => X"a88b0000",
		16#1bce# => X"8521fffc",
		16#1bcf# => X"0000012f",
		16#1bd0# => X"a8a5b838",
		16#1bd1# => X"18600001",
		16#1bd2# => X"a863b838",
		16#1bd3# => X"85630000",
		16#1bd4# => X"18600001",
		16#1bd5# => X"a863b83c",
		16#1bd6# => X"84630000",
		16#1bd7# => X"44004800",
		16#1bd8# => X"e16b1802",
		16#1bd9# => X"d7e117f8",
		16#1bda# => X"18400001",
		16#1bdb# => X"d7e14ffc",
		16#1bdc# => X"9c21fff8",
		16#1bdd# => X"0400144b",
		16#1bde# => X"a84284e8",
		16#1bdf# => X"84a20000",
		16#1be0# => X"84c20004",
		16#1be1# => X"e06b0004",
		16#1be2# => X"e08c0004",
		16#1be3# => X"04001229",
		16#1be4# => X"15000000",
		16#1be5# => X"9c210008",
		16#1be6# => X"a84b0000",
		16#1be7# => X"a86c0000",
		16#1be8# => X"8521fffc",
		16#1be9# => X"e1620004",
		16#1bea# => X"e1830004",
		16#1beb# => X"44004800",
		16#1bec# => X"8441fff8",
		16#1bed# => X"d7e117f4",
		16#1bee# => X"a8430000",
		16#1bef# => X"9c600001",
		16#1bf0# => X"d7e14ffc",
		16#1bf1# => X"d7e177f8",
		16#1bf2# => X"d8021804",
		16#1bf3# => X"040009a6",
		16#1bf4# => X"9c21fff0",
		16#1bf5# => X"18a00001",
		16#1bf6# => X"bc2b0000",
		16#1bf7# => X"0c000022",
		16#1bf8# => X"a8a5b834",
		16#1bf9# => X"84850000",
		16#1bfa# => X"bc040000",
		16#1bfb# => X"13fffffe",
		16#1bfc# => X"18800001",
		16#1bfd# => X"b9cb0002",
		16#1bfe# => X"a884b810",
		16#1bff# => X"e06e2000",
		16#1c00# => X"84a30000",
		16#1c01# => X"84850044",
		16#1c02# => X"bc240001",
		16#1c03# => X"13fffffe",
		16#1c04# => X"15000000",
		16#1c05# => X"07fff050",
		16#1c06# => X"a8650000",
		16#1c07# => X"18600001",
		16#1c08# => X"9c800000",
		16#1c09# => X"a863b810",
		16#1c0a# => X"e1ce1800",
		16#1c0b# => X"846e0000",
		16#1c0c# => X"d8022004",
		16#1c0d# => X"9c400002",
		16#1c0e# => X"d4031044",
		16#1c0f# => X"0400098a",
		16#1c10# => X"15000000",
		16#1c11# => X"bc0b0000",
		16#1c12# => X"0c000023",
		16#1c13# => X"a86b0000",
		16#1c14# => X"9c210010",
		16#1c15# => X"8521fffc",
		16#1c16# => X"8441fff4",
		16#1c17# => X"00000993",
		16#1c18# => X"85c1fff8",
		16#1c19# => X"04000980",
		16#1c1a# => X"15000000",
		16#1c1b# => X"bc0b0000",
		16#1c1c# => X"0c000013",
		16#1c1d# => X"15000000",
		16#1c1e# => X"0400097b",
		16#1c1f# => X"15000000",
		16#1c20# => X"18600001",
		16#1c21# => X"d4015800",
		16#1c22# => X"0400195c",
		16#1c23# => X"a8637ebc",
		16#1c24# => X"0400096f",
		16#1c25# => X"15000000",
		16#1c26# => X"18600001",
		16#1c27# => X"d4015800",
		16#1c28# => X"04001956",
		16#1c29# => X"a86384c0",
		16#1c2a# => X"9c210010",
		16#1c2b# => X"8521fffc",
		16#1c2c# => X"8441fff4",
		16#1c2d# => X"44004800",
		16#1c2e# => X"85c1fff8",
		16#1c2f# => X"0400096a",
		16#1c30# => X"15000000",
		16#1c31# => X"0400096e",
		16#1c32# => X"9c6bffff",
		16#1c33# => X"03ffffeb",
		16#1c34# => X"15000000",
		16#1c35# => X"0400096a",
		16#1c36# => X"9c600000",
		16#1c37# => X"0400152e",
		16#1c38# => X"9c600000",
		16#1c39# => X"d7e117f8",
		16#1c3a# => X"9c400000",
		16#1c3b# => X"d7e14ffc",
		16#1c3c# => X"d8031004",
		16#1c3d# => X"0400095c",
		16#1c3e# => X"9c21fff8",
		16#1c3f# => X"bc0b0000",
		16#1c40# => X"0c000006",
		16#1c41# => X"a86b0000",
		16#1c42# => X"9c210008",
		16#1c43# => X"8521fffc",
		16#1c44# => X"00000966",
		16#1c45# => X"8441fff8",
		16#1c46# => X"04000959",
		16#1c47# => X"9c600000",
		16#1c48# => X"0400151d",
		16#1c49# => X"9c600000",
		16#1c4a# => X"d7e117f4",
		16#1c4b# => X"18400001",
		16#1c4c# => X"d7e14ffc",
		16#1c4d# => X"a842b830",
		16#1c4e# => X"d7e177f8",
		16#1c4f# => X"84c20000",
		16#1c50# => X"bc060000",
		16#1c51# => X"10000018",
		16#1c52# => X"9c21fff4",
		16#1c53# => X"18600001",
		16#1c54# => X"a863ade0",
		16#1c55# => X"85030000",
		16#1c56# => X"19a00001",
		16#1c57# => X"b8660002",
		16#1c58# => X"a9adb810",
		16#1c59# => X"9c800001",
		16#1c5a# => X"e0636800",
		16#1c5b# => X"9d08ffff",
		16#1c5c# => X"84630000",
		16#1c5d# => X"a9cd0000",
		16#1c5e# => X"d4032044",
		16#1c5f# => X"e4264000",
		16#1c60# => X"0c000025",
		16#1c61# => X"9cc60001",
		16#1c62# => X"9d600000",
		16#1c63# => X"d4023000",
		16#1c64# => X"9c21000c",
		16#1c65# => X"8521fffc",
		16#1c66# => X"8441fff4",
		16#1c67# => X"44004800",
		16#1c68# => X"85c1fff8",
		16#1c69# => X"18800001",
		16#1c6a# => X"a884ade0",
		16#1c6b# => X"85040000",
		16#1c6c# => X"bc080000",
		16#1c6d# => X"10000012",
		16#1c6e# => X"a8860000",
		16#1c6f# => X"a8a60000",
		16#1c70# => X"9d80004c",
		16#1c71# => X"e0e56306",
		16#1c72# => X"19a00001",
		16#1c73# => X"b8a50002",
		16#1c74# => X"a9adb810",
		16#1c75# => X"e0e33800",
		16#1c76# => X"e1656800",
		16#1c77# => X"9c840001",
		16#1c78# => X"d40b3800",
		16#1c79# => X"9d600000",
		16#1c7a# => X"a8a40000",
		16#1c7b# => X"d4075844",
		16#1c7c# => X"e4244000",
		16#1c7d# => X"13fffff5",
		16#1c7e# => X"e0e56306",
		16#1c7f# => X"18600001",
		16#1c80# => X"9c800001",
		16#1c81# => X"a863b834",
		16#1c82# => X"d4032000",
		16#1c83# => X"03ffffd4",
		16#1c84# => X"19a00001",
		16#1c85# => X"07ffefd0",
		16#1c86# => X"846d0000",
		16#1c87# => X"84c20000",
		16#1c88# => X"846e0000",
		16#1c89# => X"9c800002",
		16#1c8a# => X"9cc60001",
		16#1c8b# => X"d4032044",
		16#1c8c# => X"d4023000",
		16#1c8d# => X"9c21000c",
		16#1c8e# => X"9d600000",
		16#1c8f# => X"8521fffc",
		16#1c90# => X"8441fff4",
		16#1c91# => X"44004800",
		16#1c92# => X"85c1fff8",
		16#1c93# => X"18a00001",
		16#1c94# => X"d7e117fc",
		16#1c95# => X"a8a5b80c",
		16#1c96# => X"18400001",
		16#1c97# => X"84c50000",
		16#1c98# => X"a842b810",
		16#1c99# => X"b8660002",
		16#1c9a# => X"9c21fffc",
		16#1c9b# => X"e0631000",
		16#1c9c# => X"84830000",
		16#1c9d# => X"84640044",
		16#1c9e# => X"bc230002",
		16#1c9f# => X"13fffffe",
		16#1ca0# => X"9d600000",
		16#1ca1# => X"9cc60001",
		16#1ca2# => X"d4053000",
		16#1ca3# => X"9c210004",
		16#1ca4# => X"44004800",
		16#1ca5# => X"8441fffc",
		16#1ca6# => X"18800001",
		16#1ca7# => X"a884b8c0",
		16#1ca8# => X"44004800",
		16#1ca9# => X"d4041800",
		16#1caa# => X"b8840004",
		16#1cab# => X"e0641800",
		16#1cac# => X"9c800001",
		16#1cad# => X"d4032000",
		16#1cae# => X"44004800",
		16#1caf# => X"15000000",
		16#1cb0# => X"b8840004",
		16#1cb1# => X"e0641800",
		16#1cb2# => X"9c800002",
		16#1cb3# => X"d4032000",
		16#1cb4# => X"44004800",
		16#1cb5# => X"15000000",
		16#1cb6# => X"b8840004",
		16#1cb7# => X"d7e117fc",
		16#1cb8# => X"9c400000",
		16#1cb9# => X"e0641800",
		16#1cba# => X"9c21fffc",
		16#1cbb# => X"d4031000",
		16#1cbc# => X"9c210004",
		16#1cbd# => X"44004800",
		16#1cbe# => X"8441fffc",
		16#1cbf# => X"b8840004",
		16#1cc0# => X"e0632000",
		16#1cc1# => X"85630004",
		16#1cc2# => X"44004800",
		16#1cc3# => X"15000000",
		16#1cc4# => X"b8c40004",
		16#1cc5# => X"9c630004",
		16#1cc6# => X"d7e117fc",
		16#1cc7# => X"e0633000",
		16#1cc8# => X"9c21fffc",
		16#1cc9# => X"d4032800",
		16#1cca# => X"9d60ffff",
		16#1ccb# => X"84630000",
		16#1ccc# => X"e4232800",
		16#1ccd# => X"10000007",
		16#1cce# => X"b8840002",
		16#1ccf# => X"18400001",
		16#1cd0# => X"a842b840",
		16#1cd1# => X"9d600000",
		16#1cd2# => X"e0841000",
		16#1cd3# => X"d4041800",
		16#1cd4# => X"9c210004",
		16#1cd5# => X"44004800",
		16#1cd6# => X"8441fffc",
		16#1cd7# => X"b8840004",
		16#1cd8# => X"e0632000",
		16#1cd9# => X"85630008",
		16#1cda# => X"44004800",
		16#1cdb# => X"15000000",
		16#1cdc# => X"18a00001",
		16#1cdd# => X"d7e117f4",
		16#1cde# => X"b8440002",
		16#1cdf# => X"a8a5b840",
		16#1ce0# => X"d7e14ffc",
		16#1ce1# => X"e0422800",
		16#1ce2# => X"d7e177f8",
		16#1ce3# => X"84420000",
		16#1ce4# => X"bc020000",
		16#1ce5# => X"0c000003",
		16#1ce6# => X"9c21fff4",
		16#1ce7# => X"9c400001",
		16#1ce8# => X"b8a40004",
		16#1ce9# => X"9c8003e8",
		16#1cea# => X"e0a32800",
		16#1ceb# => X"18600001",
		16#1cec# => X"85c50008",
		16#1ced# => X"a863b8c0",
		16#1cee# => X"0400091d",
		16#1cef# => X"84630000",
		16#1cf0# => X"a86e0000",
		16#1cf1# => X"040008db",
		16#1cf2# => X"a88b0000",
		16#1cf3# => X"9c21000c",
		16#1cf4# => X"e1625b06",
		16#1cf5# => X"8521fffc",
		16#1cf6# => X"8441fff4",
		16#1cf7# => X"44004800",
		16#1cf8# => X"85c1fff8",
		16#1cf9# => X"b8840004",
		16#1cfa# => X"e0632000",
		16#1cfb# => X"84630008",
		16#1cfc# => X"44004800",
		16#1cfd# => X"d4051800",
		16#1cfe# => X"d7e177f4",
		16#1cff# => X"a9c50000",
		16#1d00# => X"18a00001",
		16#1d01# => X"d7e117f0",
		16#1d02# => X"b8440002",
		16#1d03# => X"a8a5b840",
		16#1d04# => X"d7e14ffc",
		16#1d05# => X"e0422800",
		16#1d06# => X"d7e187f8",
		16#1d07# => X"84420000",
		16#1d08# => X"bc020000",
		16#1d09# => X"0c000003",
		16#1d0a# => X"9c21fff0",
		16#1d0b# => X"9c400001",
		16#1d0c# => X"b8a40004",
		16#1d0d# => X"9c8003e8",
		16#1d0e# => X"e0a32800",
		16#1d0f# => X"18600001",
		16#1d10# => X"86050008",
		16#1d11# => X"a863b8c0",
		16#1d12# => X"040008f9",
		16#1d13# => X"84630000",
		16#1d14# => X"a8700000",
		16#1d15# => X"040008b7",
		16#1d16# => X"a88b0000",
		16#1d17# => X"e0425b06",
		16#1d18# => X"d40e1000",
		16#1d19# => X"9c210010",
		16#1d1a# => X"8521fffc",
		16#1d1b# => X"8441fff0",
		16#1d1c# => X"85c1fff4",
		16#1d1d# => X"44004800",
		16#1d1e# => X"8601fff8",
		16#1d1f# => X"d7e14ffc",
		16#1d20# => X"9c21fffc",
		16#1d21# => X"a860c800",
		16#1d22# => X"9c210004",
		16#1d23# => X"8521fffc",
		16#1d24# => X"000017f4",
		16#1d25# => X"9c800001",
		16#1d26# => X"d7e14ffc",
		16#1d27# => X"9c21fffc",
		16#1d28# => X"a860c800",
		16#1d29# => X"9c210004",
		16#1d2a# => X"8521fffc",
		16#1d2b# => X"000017ed",
		16#1d2c# => X"9c800000",
		16#1d2d# => X"d7e177f8",
		16#1d2e# => X"a9c40000",
		16#1d2f# => X"a880c83e",
		16#1d30# => X"d7e14ffc",
		16#1d31# => X"d7e117f4",
		16#1d32# => X"9c21fff4",
		16#1d33# => X"a8430000",
		16#1d34# => X"040017e7",
		16#1d35# => X"e06e2000",
		16#1d36# => X"a880c83c",
		16#1d37# => X"d4025800",
		16#1d38# => X"040017e3",
		16#1d39# => X"e06e2000",
		16#1d3a# => X"a880c83d",
		16#1d3b# => X"9d6b0001",
		16#1d3c# => X"e06e2000",
		16#1d3d# => X"040017de",
		16#1d3e# => X"d4025804",
		16#1d3f# => X"a880c83f",
		16#1d40# => X"9d6b0001",
		16#1d41# => X"e06e2000",
		16#1d42# => X"040017d9",
		16#1d43# => X"d402580c",
		16#1d44# => X"a86b0000",
		16#1d45# => X"04000cb6",
		16#1d46# => X"d4025810",
		16#1d47# => X"84620000",
		16#1d48# => X"04000cb3",
		16#1d49# => X"a9cb0000",
		16#1d4a# => X"a86e0000",
		16#1d4b# => X"04000b05",
		16#1d4c# => X"a88b0000",
		16#1d4d# => X"d4025808",
		16#1d4e# => X"9c21000c",
		16#1d4f# => X"8521fffc",
		16#1d50# => X"8441fff4",
		16#1d51# => X"44004800",
		16#1d52# => X"85c1fff8",
		16#1d53# => X"d7e14ffc",
		16#1d54# => X"d7e117d4",
		16#1d55# => X"d7e177d8",
		16#1d56# => X"d7e187dc",
		16#1d57# => X"d7e197e0",
		16#1d58# => X"d7e1a7e4",
		16#1d59# => X"d7e1b7e8",
		16#1d5a# => X"d7e1c7ec",
		16#1d5b# => X"d7e1d7f0",
		16#1d5c# => X"d7e1e7f4",
		16#1d5d# => X"d7e1f7f8",
		16#1d5e# => X"0400083b",
		16#1d5f# => X"9c21ff74",
		16#1d60# => X"a860c87e",
		16#1d61# => X"040017ba",
		16#1d62# => X"a84b0000",
		16#1d63# => X"b8820002",
		16#1d64# => X"b8420004",
		16#1d65# => X"a860c87c",
		16#1d66# => X"e2c41000",
		16#1d67# => X"18400001",
		16#1d68# => X"18800001",
		16#1d69# => X"a842b8c4",
		16#1d6a# => X"a884ba2c",
		16#1d6b# => X"e0561000",
		16#1d6c# => X"e0962000",
		16#1d6d# => X"d4025800",
		16#1d6e# => X"d4012004",
		16#1d6f# => X"040017ac",
		16#1d70# => X"d4011000",
		16#1d71# => X"9d6b0001",
		16#1d72# => X"a860c87d",
		16#1d73# => X"9ca20010",
		16#1d74# => X"d4025804",
		16#1d75# => X"040017a6",
		16#1d76# => X"d4012824",
		16#1d77# => X"9d6b0001",
		16#1d78# => X"a860c87f",
		16#1d79# => X"d402580c",
		16#1d7a# => X"040017a1",
		16#1d7b# => X"9e020008",
		16#1d7c# => X"84c10004",
		16#1d7d# => X"84410024",
		16#1d7e# => X"9cc60010",
		16#1d7f# => X"a86b0000",
		16#1d80# => X"d4025800",
		16#1d81# => X"04000c7a",
		16#1d82# => X"d4013028",
		16#1d83# => X"84810000",
		16#1d84# => X"84a10004",
		16#1d85# => X"84640000",
		16#1d86# => X"9dc50008",
		16#1d87# => X"04000c74",
		16#1d88# => X"aa4b0000",
		16#1d89# => X"18c00001",
		16#1d8a# => X"a88b0000",
		16#1d8b# => X"a8c6bae0",
		16#1d8c# => X"a8720000",
		16#1d8d# => X"04000ac3",
		16#1d8e# => X"e3d63000",
		16#1d8f# => X"a860c8be",
		16#1d90# => X"d4105800",
		16#1d91# => X"0400178a",
		16#1d92# => X"9e5e0008",
		16#1d93# => X"84410004",
		16#1d94# => X"a860c8bc",
		16#1d95# => X"04001786",
		16#1d96# => X"d4025800",
		16#1d97# => X"9d6b0001",
		16#1d98# => X"a860c8bd",
		16#1d99# => X"9c9e0010",
		16#1d9a# => X"d4025804",
		16#1d9b# => X"04001780",
		16#1d9c# => X"d401202c",
		16#1d9d# => X"9d6b0001",
		16#1d9e# => X"a860c8bf",
		16#1d9f# => X"0400177c",
		16#1da0# => X"d402580c",
		16#1da1# => X"18a00001",
		16#1da2# => X"84c10028",
		16#1da3# => X"a8a5bb94",
		16#1da4# => X"d4065800",
		16#1da5# => X"a86b0000",
		16#1da6# => X"04000c55",
		16#1da7# => X"e3962800",
		16#1da8# => X"84620000",
		16#1da9# => X"9c5c0010",
		16#1daa# => X"aa0b0000",
		16#1dab# => X"04000c50",
		16#1dac# => X"d4011030",
		16#1dad# => X"a8700000",
		16#1dae# => X"a88b0000",
		16#1daf# => X"04000aa1",
		16#1db0# => X"18400001",
		16#1db1# => X"a860c8fe",
		16#1db2# => X"d40e5800",
		16#1db3# => X"04001768",
		16#1db4# => X"a842bcfc",
		16#1db5# => X"a860c8fc",
		16#1db6# => X"d41e5800",
		16#1db7# => X"04001764",
		16#1db8# => X"e3161000",
		16#1db9# => X"18800001",
		16#1dba# => X"9d6b0001",
		16#1dbb# => X"a860c8fd",
		16#1dbc# => X"a884bc48",
		16#1dbd# => X"d41e5804",
		16#1dbe# => X"0400175d",
		16#1dbf# => X"e3562000",
		16#1dc0# => X"9d6b0001",
		16#1dc1# => X"a860c8ff",
		16#1dc2# => X"9cba0010",
		16#1dc3# => X"d41e580c",
		16#1dc4# => X"04001757",
		16#1dc5# => X"d4012834",
		16#1dc6# => X"84c1002c",
		16#1dc7# => X"a86b0000",
		16#1dc8# => X"d4065800",
		16#1dc9# => X"04000c32",
		16#1dca# => X"9e1c0008",
		16#1dcb# => X"847e0000",
		16#1dcc# => X"04000c2f",
		16#1dcd# => X"aa8b0000",
		16#1dce# => X"9cb80010",
		16#1dcf# => X"a88b0000",
		16#1dd0# => X"a8740000",
		16#1dd1# => X"04000a7f",
		16#1dd2# => X"d4012838",
		16#1dd3# => X"a860c93e",
		16#1dd4# => X"d4125800",
		16#1dd5# => X"04001746",
		16#1dd6# => X"9dda0008",
		16#1dd7# => X"a860c93c",
		16#1dd8# => X"d41c5800",
		16#1dd9# => X"04001742",
		16#1dda# => X"9c580008",
		16#1ddb# => X"9d6b0001",
		16#1ddc# => X"a860c93d",
		16#1ddd# => X"0400173e",
		16#1dde# => X"d41c5804",
		16#1ddf# => X"18c00001",
		16#1de0# => X"9d6b0001",
		16#1de1# => X"a8c6bdb0",
		16#1de2# => X"a860c93f",
		16#1de3# => X"d41c580c",
		16#1de4# => X"04001737",
		16#1de5# => X"e2963000",
		16#1de6# => X"84810030",
		16#1de7# => X"9c740010",
		16#1de8# => X"d4045800",
		16#1de9# => X"d401183c",
		16#1dea# => X"04000c11",
		16#1deb# => X"a86b0000",
		16#1dec# => X"9cb40008",
		16#1ded# => X"847c0000",
		16#1dee# => X"d4012820",
		16#1def# => X"04000c0c",
		16#1df0# => X"aa4b0000",
		16#1df1# => X"18c00001",
		16#1df2# => X"a88b0000",
		16#1df3# => X"a8c6be64",
		16#1df4# => X"a8720000",
		16#1df5# => X"04000a5b",
		16#1df6# => X"e2563000",
		16#1df7# => X"a860c97e",
		16#1df8# => X"04001723",
		16#1df9# => X"d4105800",
		16#1dfa# => X"a860c97c",
		16#1dfb# => X"04001720",
		16#1dfc# => X"d41a5800",
		16#1dfd# => X"9d6b0001",
		16#1dfe# => X"a860c97d",
		16#1dff# => X"9c920008",
		16#1e00# => X"d41a5804",
		16#1e01# => X"0400171a",
		16#1e02# => X"d4012040",
		16#1e03# => X"18a00001",
		16#1e04# => X"9d6b0001",
		16#1e05# => X"a8a5c350",
		16#1e06# => X"a860c97f",
		16#1e07# => X"e0b62800",
		16#1e08# => X"d41a580c",
		16#1e09# => X"04001712",
		16#1e0a# => X"d4012808",
		16#1e0b# => X"84810034",
		16#1e0c# => X"84c10008",
		16#1e0d# => X"d4045800",
		16#1e0e# => X"9cc60008",
		16#1e0f# => X"a86b0000",
		16#1e10# => X"04000beb",
		16#1e11# => X"d4013044",
		16#1e12# => X"18a00001",
		16#1e13# => X"847a0000",
		16#1e14# => X"a8a5c404",
		16#1e15# => X"aa0b0000",
		16#1e16# => X"e0b62800",
		16#1e17# => X"04000be4",
		16#1e18# => X"d401280c",
		16#1e19# => X"84c1000c",
		16#1e1a# => X"a88b0000",
		16#1e1b# => X"9cc60008",
		16#1e1c# => X"a8700000",
		16#1e1d# => X"04000a33",
		16#1e1e# => X"d4013048",
		16#1e1f# => X"a860c9be",
		16#1e20# => X"040016fb",
		16#1e21# => X"d40e5800",
		16#1e22# => X"a860c9bc",
		16#1e23# => X"040016f8",
		16#1e24# => X"d4185800",
		16#1e25# => X"18800001",
		16#1e26# => X"9d6b0001",
		16#1e27# => X"a884bf18",
		16#1e28# => X"a860c9bd",
		16#1e29# => X"e0962000",
		16#1e2a# => X"d4185804",
		16#1e2b# => X"040016f0",
		16#1e2c# => X"d4012010",
		16#1e2d# => X"84a10010",
		16#1e2e# => X"9d6b0001",
		16#1e2f# => X"a860c9bf",
		16#1e30# => X"9ca50008",
		16#1e31# => X"d418580c",
		16#1e32# => X"040016e9",
		16#1e33# => X"d401284c",
		16#1e34# => X"18c00001",
		16#1e35# => X"84810038",
		16#1e36# => X"a8c6bfcc",
		16#1e37# => X"d4045800",
		16#1e38# => X"e0d63000",
		16#1e39# => X"a86b0000",
		16#1e3a# => X"04000bc1",
		16#1e3b# => X"d4013014",
		16#1e3c# => X"84a10014",
		16#1e3d# => X"84780000",
		16#1e3e# => X"9ca50008",
		16#1e3f# => X"a9cb0000",
		16#1e40# => X"04000bbb",
		16#1e41# => X"d4012850",
		16#1e42# => X"18c00001",
		16#1e43# => X"a88b0000",
		16#1e44# => X"a8c6c080",
		16#1e45# => X"a86e0000",
		16#1e46# => X"e0d63000",
		16#1e47# => X"04000a09",
		16#1e48# => X"d4013018",
		16#1e49# => X"a860c9fe",
		16#1e4a# => X"040016d1",
		16#1e4b# => X"d4025800",
		16#1e4c# => X"a860c9fc",
		16#1e4d# => X"040016ce",
		16#1e4e# => X"d4145800",
		16#1e4f# => X"84410018",
		16#1e50# => X"9d6b0001",
		16#1e51# => X"a860c9fd",
		16#1e52# => X"9c420008",
		16#1e53# => X"d4145804",
		16#1e54# => X"040016c7",
		16#1e55# => X"d4011054",
		16#1e56# => X"18800001",
		16#1e57# => X"9d6b0001",
		16#1e58# => X"a884c134",
		16#1e59# => X"a860c9ff",
		16#1e5a# => X"e0962000",
		16#1e5b# => X"d414580c",
		16#1e5c# => X"040016bf",
		16#1e5d# => X"d401201c",
		16#1e5e# => X"84c1003c",
		16#1e5f# => X"84a1001c",
		16#1e60# => X"d4065800",
		16#1e61# => X"9ca50008",
		16#1e62# => X"a86b0000",
		16#1e63# => X"18400001",
		16#1e64# => X"d4012858",
		16#1e65# => X"04000b96",
		16#1e66# => X"a842c1e8",
		16#1e67# => X"84740000",
		16#1e68# => X"e2161000",
		16#1e69# => X"04000b92",
		16#1e6a# => X"a9cb0000",
		16#1e6b# => X"9cb00008",
		16#1e6c# => X"a88b0000",
		16#1e6d# => X"a86e0000",
		16#1e6e# => X"040009e2",
		16#1e6f# => X"d401285c",
		16#1e70# => X"84c10020",
		16#1e71# => X"a860ca3e",
		16#1e72# => X"040016a9",
		16#1e73# => X"d4065800",
		16#1e74# => X"a860ca3c",
		16#1e75# => X"040016a6",
		16#1e76# => X"d4125800",
		16#1e77# => X"18800001",
		16#1e78# => X"9d6b0001",
		16#1e79# => X"a860ca3d",
		16#1e7a# => X"a884c29c",
		16#1e7b# => X"d4125804",
		16#1e7c# => X"0400169f",
		16#1e7d# => X"e0562000",
		16#1e7e# => X"9d6b0001",
		16#1e7f# => X"a860ca3f",
		16#1e80# => X"9ca20008",
		16#1e81# => X"d412580c",
		16#1e82# => X"04001699",
		16#1e83# => X"d4012820",
		16#1e84# => X"a86b0000",
		16#1e85# => X"04000b76",
		16#1e86# => X"d4125810",
		16#1e87# => X"84720000",
		16#1e88# => X"04000b73",
		16#1e89# => X"a9cb0000",
		16#1e8a# => X"a86e0000",
		16#1e8b# => X"040009c5",
		16#1e8c# => X"a88b0000",
		16#1e8d# => X"84c10040",
		16#1e8e# => X"a860ca7e",
		16#1e8f# => X"0400168c",
		16#1e90# => X"d4065800",
		16#1e91# => X"84810008",
		16#1e92# => X"a860ca7c",
		16#1e93# => X"04001688",
		16#1e94# => X"d4045800",
		16#1e95# => X"84a10008",
		16#1e96# => X"9d6b0001",
		16#1e97# => X"a860ca7d",
		16#1e98# => X"04001683",
		16#1e99# => X"d4055804",
		16#1e9a# => X"84c10008",
		16#1e9b# => X"9d6b0001",
		16#1e9c# => X"a860ca7f",
		16#1e9d# => X"0400167e",
		16#1e9e# => X"d406580c",
		16#1e9f# => X"84810008",
		16#1ea0# => X"a86b0000",
		16#1ea1# => X"04000b5a",
		16#1ea2# => X"d4045810",
		16#1ea3# => X"84a10008",
		16#1ea4# => X"a9cb0000",
		16#1ea5# => X"04000b56",
		16#1ea6# => X"84650000",
		16#1ea7# => X"a86e0000",
		16#1ea8# => X"040009a8",
		16#1ea9# => X"a88b0000",
		16#1eaa# => X"84c10044",
		16#1eab# => X"a860cabe",
		16#1eac# => X"0400166f",
		16#1ead# => X"d4065800",
		16#1eae# => X"8481000c",
		16#1eaf# => X"a860cabc",
		16#1eb0# => X"0400166b",
		16#1eb1# => X"d4045800",
		16#1eb2# => X"84a1000c",
		16#1eb3# => X"9d6b0001",
		16#1eb4# => X"a860cabd",
		16#1eb5# => X"04001666",
		16#1eb6# => X"d4055804",
		16#1eb7# => X"84c1000c",
		16#1eb8# => X"9d6b0001",
		16#1eb9# => X"a860cabf",
		16#1eba# => X"04001661",
		16#1ebb# => X"d406580c",
		16#1ebc# => X"8481000c",
		16#1ebd# => X"a86b0000",
		16#1ebe# => X"04000b3d",
		16#1ebf# => X"d4045810",
		16#1ec0# => X"84a1000c",
		16#1ec1# => X"a9cb0000",
		16#1ec2# => X"04000b39",
		16#1ec3# => X"84650000",
		16#1ec4# => X"a86e0000",
		16#1ec5# => X"0400098b",
		16#1ec6# => X"a88b0000",
		16#1ec7# => X"84c10048",
		16#1ec8# => X"a860cafe",
		16#1ec9# => X"04001652",
		16#1eca# => X"d4065800",
		16#1ecb# => X"84810010",
		16#1ecc# => X"a860cafc",
		16#1ecd# => X"0400164e",
		16#1ece# => X"d4045800",
		16#1ecf# => X"84a10010",
		16#1ed0# => X"9d6b0001",
		16#1ed1# => X"a860cafd",
		16#1ed2# => X"04001649",
		16#1ed3# => X"d4055804",
		16#1ed4# => X"84c10010",
		16#1ed5# => X"9d6b0001",
		16#1ed6# => X"a860caff",
		16#1ed7# => X"04001644",
		16#1ed8# => X"d406580c",
		16#1ed9# => X"84810010",
		16#1eda# => X"a86b0000",
		16#1edb# => X"04000b20",
		16#1edc# => X"d4045810",
		16#1edd# => X"84a10010",
		16#1ede# => X"a9cb0000",
		16#1edf# => X"04000b1c",
		16#1ee0# => X"84650000",
		16#1ee1# => X"a86e0000",
		16#1ee2# => X"0400096e",
		16#1ee3# => X"a88b0000",
		16#1ee4# => X"84c1004c",
		16#1ee5# => X"a860cb3e",
		16#1ee6# => X"04001635",
		16#1ee7# => X"d4065800",
		16#1ee8# => X"84810014",
		16#1ee9# => X"a860cb3c",
		16#1eea# => X"04001631",
		16#1eeb# => X"d4045800",
		16#1eec# => X"84a10014",
		16#1eed# => X"9d6b0001",
		16#1eee# => X"a860cb3d",
		16#1eef# => X"0400162c",
		16#1ef0# => X"d4055804",
		16#1ef1# => X"84c10014",
		16#1ef2# => X"9d6b0001",
		16#1ef3# => X"a860cb3f",
		16#1ef4# => X"04001627",
		16#1ef5# => X"d406580c",
		16#1ef6# => X"84810014",
		16#1ef7# => X"a86b0000",
		16#1ef8# => X"04000b03",
		16#1ef9# => X"d4045810",
		16#1efa# => X"84a10014",
		16#1efb# => X"a9cb0000",
		16#1efc# => X"04000aff",
		16#1efd# => X"84650000",
		16#1efe# => X"a86e0000",
		16#1eff# => X"04000951",
		16#1f00# => X"a88b0000",
		16#1f01# => X"84c10050",
		16#1f02# => X"a860cb7e",
		16#1f03# => X"04001618",
		16#1f04# => X"d4065800",
		16#1f05# => X"84810018",
		16#1f06# => X"a860cb7c",
		16#1f07# => X"04001614",
		16#1f08# => X"d4045800",
		16#1f09# => X"84a10018",
		16#1f0a# => X"9d6b0001",
		16#1f0b# => X"a860cb7d",
		16#1f0c# => X"0400160f",
		16#1f0d# => X"d4055804",
		16#1f0e# => X"84c10018",
		16#1f0f# => X"9d6b0001",
		16#1f10# => X"a860cb7f",
		16#1f11# => X"0400160a",
		16#1f12# => X"d406580c",
		16#1f13# => X"84810018",
		16#1f14# => X"a86b0000",
		16#1f15# => X"04000ae6",
		16#1f16# => X"d4045810",
		16#1f17# => X"84a10018",
		16#1f18# => X"a9cb0000",
		16#1f19# => X"04000ae2",
		16#1f1a# => X"84650000",
		16#1f1b# => X"a86e0000",
		16#1f1c# => X"04000934",
		16#1f1d# => X"a88b0000",
		16#1f1e# => X"84c10054",
		16#1f1f# => X"a860cbbe",
		16#1f20# => X"040015fb",
		16#1f21# => X"d4065800",
		16#1f22# => X"8481001c",
		16#1f23# => X"a860cbbc",
		16#1f24# => X"040015f7",
		16#1f25# => X"d4045800",
		16#1f26# => X"84a1001c",
		16#1f27# => X"9d6b0001",
		16#1f28# => X"a860cbbd",
		16#1f29# => X"040015f2",
		16#1f2a# => X"d4055804",
		16#1f2b# => X"84c1001c",
		16#1f2c# => X"9d6b0001",
		16#1f2d# => X"a860cbbf",
		16#1f2e# => X"040015ed",
		16#1f2f# => X"d406580c",
		16#1f30# => X"8481001c",
		16#1f31# => X"a86b0000",
		16#1f32# => X"04000ac9",
		16#1f33# => X"d4045810",
		16#1f34# => X"84a1001c",
		16#1f35# => X"a9cb0000",
		16#1f36# => X"04000ac5",
		16#1f37# => X"84650000",
		16#1f38# => X"a86e0000",
		16#1f39# => X"04000917",
		16#1f3a# => X"a88b0000",
		16#1f3b# => X"84c10058",
		16#1f3c# => X"a860cbfe",
		16#1f3d# => X"040015de",
		16#1f3e# => X"d4065800",
		16#1f3f# => X"a860cbfc",
		16#1f40# => X"040015db",
		16#1f41# => X"d4105800",
		16#1f42# => X"9d6b0001",
		16#1f43# => X"a860cbfd",
		16#1f44# => X"040015d7",
		16#1f45# => X"d4105804",
		16#1f46# => X"9d6b0001",
		16#1f47# => X"a860cbff",
		16#1f48# => X"040015d3",
		16#1f49# => X"d410580c",
		16#1f4a# => X"a86b0000",
		16#1f4b# => X"04000ab0",
		16#1f4c# => X"d4105810",
		16#1f4d# => X"84700000",
		16#1f4e# => X"04000aad",
		16#1f4f# => X"a9cb0000",
		16#1f50# => X"a86e0000",
		16#1f51# => X"040008ff",
		16#1f52# => X"a88b0000",
		16#1f53# => X"8481005c",
		16#1f54# => X"a860cc3e",
		16#1f55# => X"040015c6",
		16#1f56# => X"d4045800",
		16#1f57# => X"a860cc3c",
		16#1f58# => X"040015c3",
		16#1f59# => X"d4025800",
		16#1f5a# => X"9d6b0001",
		16#1f5b# => X"a860cc3d",
		16#1f5c# => X"040015bf",
		16#1f5d# => X"d4025804",
		16#1f5e# => X"9d6b0001",
		16#1f5f# => X"a860cc3f",
		16#1f60# => X"040015bb",
		16#1f61# => X"d402580c",
		16#1f62# => X"a86b0000",
		16#1f63# => X"04000a98",
		16#1f64# => X"d4025810",
		16#1f65# => X"84620000",
		16#1f66# => X"04000a95",
		16#1f67# => X"a9cb0000",
		16#1f68# => X"a86e0000",
		16#1f69# => X"040008e7",
		16#1f6a# => X"a88b0000",
		16#1f6b# => X"84c10028",
		16#1f6c# => X"84410024",
		16#1f6d# => X"84a60000",
		16#1f6e# => X"84620000",
		16#1f6f# => X"8481002c",
		16#1f70# => X"e0a51800",
		16#1f71# => X"84c40000",
		16#1f72# => X"84610004",
		16#1f73# => X"84810000",
		16#1f74# => X"84430000",
		16#1f75# => X"84640000",
		16#1f76# => X"e0a53000",
		16#1f77# => X"e0421800",
		16#1f78# => X"84610030",
		16#1f79# => X"84810034",
		16#1f7a# => X"84c30000",
		16#1f7b# => X"847e0000",
		16#1f7c# => X"e0a53000",
		16#1f7d# => X"e0421800",
		16#1f7e# => X"847c0000",
		16#1f7f# => X"84c40000",
		16#1f80# => X"e0421800",
		16#1f81# => X"84610038",
		16#1f82# => X"8481003c",
		16#1f83# => X"e0a53000",
		16#1f84# => X"84c30000",
		16#1f85# => X"847a0000",
		16#1f86# => X"e0a53000",
		16#1f87# => X"84c40000",
		16#1f88# => X"e0421800",
		16#1f89# => X"e0a53000",
		16#1f8a# => X"84780000",
		16#1f8b# => X"18c00001",
		16#1f8c# => X"e0421800",
		16#1f8d# => X"a8c6b978",
		16#1f8e# => X"84740000",
		16#1f8f# => X"e0963000",
		16#1f90# => X"e0421800",
		16#1f91# => X"84c10020",
		16#1f92# => X"a8650000",
		16#1f93# => X"d4042810",
		16#1f94# => X"d4041000",
		16#1f95# => X"d4065800",
		16#1f96# => X"04000a65",
		16#1f97# => X"9dc40008",
		16#1f98# => X"a8620000",
		16#1f99# => X"04000a62",
		16#1f9a# => X"aa0b0000",
		16#1f9b# => X"a8700000",
		16#1f9c# => X"040008b4",
		16#1f9d# => X"a88b0000",
		16#1f9e# => X"d40e5800",
		16#1f9f# => X"9c21008c",
		16#1fa0# => X"8521fffc",
		16#1fa1# => X"8441ffd4",
		16#1fa2# => X"85c1ffd8",
		16#1fa3# => X"8601ffdc",
		16#1fa4# => X"8641ffe0",
		16#1fa5# => X"8681ffe4",
		16#1fa6# => X"86c1ffe8",
		16#1fa7# => X"8701ffec",
		16#1fa8# => X"8741fff0",
		16#1fa9# => X"8781fff4",
		16#1faa# => X"44004800",
		16#1fab# => X"87c1fff8",
		16#1fac# => X"d7e14ffc",
		16#1fad# => X"d7e117d4",
		16#1fae# => X"d7e177d8",
		16#1faf# => X"d7e187dc",
		16#1fb0# => X"d7e197e0",
		16#1fb1# => X"d7e1a7e4",
		16#1fb2# => X"d7e1b7e8",
		16#1fb3# => X"d7e1c7ec",
		16#1fb4# => X"d7e1d7f0",
		16#1fb5# => X"d7e1e7f4",
		16#1fb6# => X"d7e1f7f8",
		16#1fb7# => X"040005e2",
		16#1fb8# => X"9c21ff98",
		16#1fb9# => X"18600001",
		16#1fba# => X"a84b0000",
		16#1fbb# => X"a86384f0",
		16#1fbc# => X"040015c2",
		16#1fbd# => X"d4015800",
		16#1fbe# => X"18600001",
		16#1fbf# => X"d4011000",
		16#1fc0# => X"a863853c",
		16#1fc1# => X"040015bd",
		16#1fc2# => X"b9c20002",
		16#1fc3# => X"18800001",
		16#1fc4# => X"18600001",
		16#1fc5# => X"a8848586",
		16#1fc6# => X"a8638560",
		16#1fc7# => X"d4012004",
		16#1fc8# => X"18800001",
		16#1fc9# => X"d4011000",
		16#1fca# => X"a884858c",
		16#1fcb# => X"d4012008",
		16#1fcc# => X"18800001",
		16#1fcd# => X"a8848592",
		16#1fce# => X"d401200c",
		16#1fcf# => X"18800001",
		16#1fd0# => X"a8848596",
		16#1fd1# => X"d4012010",
		16#1fd2# => X"18800001",
		16#1fd3# => X"a884859a",
		16#1fd4# => X"d4012014",
		16#1fd5# => X"18800001",
		16#1fd6# => X"a884859e",
		16#1fd7# => X"d4012018",
		16#1fd8# => X"18800001",
		16#1fd9# => X"a88485a4",
		16#1fda# => X"040015a4",
		16#1fdb# => X"d401201c",
		16#1fdc# => X"18600001",
		16#1fdd# => X"d4011000",
		16#1fde# => X"040015a0",
		16#1fdf# => X"a86384f0",
		16#1fe0# => X"b8620004",
		16#1fe1# => X"18800001",
		16#1fe2# => X"d4011000",
		16#1fe3# => X"e1ce1800",
		16#1fe4# => X"18600001",
		16#1fe5# => X"a884b978",
		16#1fe6# => X"a86385d3",
		16#1fe7# => X"e08e2000",
		16#1fe8# => X"d4011804",
		16#1fe9# => X"18600001",
		16#1fea# => X"d4012030",
		16#1feb# => X"a863b8c4",
		16#1fec# => X"e20e1800",
		16#1fed# => X"84700008",
		16#1fee# => X"84b00000",
		16#1fef# => X"84900004",
		16#1ff0# => X"86500010",
		16#1ff1# => X"d4012808",
		16#1ff2# => X"04000a96",
		16#1ff3# => X"d401200c",
		16#1ff4# => X"8490000c",
		16#1ff5# => X"84a10030",
		16#1ff6# => X"a8720000",
		16#1ff7# => X"9ec50010",
		16#1ff8# => X"d4015810",
		16#1ff9# => X"d4016014",
		16#1ffa# => X"d4012018",
		16#1ffb# => X"04000a00",
		16#1ffc# => X"d401901c",
		16#1ffd# => X"18c00001",
		16#1ffe# => X"84760000",
		16#1fff# => X"a8c6ba2c",
		16#2000# => X"aa4b0000",
		16#2001# => X"040009fa",
		16#2002# => X"e20e3000",
		16#2003# => X"18a00001",
		16#2004# => X"a88b0000",
		16#2005# => X"a8a5bae0",
		16#2006# => X"a8720000",
		16#2007# => X"04000849",
		16#2008# => X"e28e2800",
		16#2009# => X"18c00001",
		16#200a# => X"a86b0000",
		16#200b# => X"a8c6bb94",
		16#200c# => X"04000a7c",
		16#200d# => X"e24e3000",
		16#200e# => X"18600001",
		16#200f# => X"d4015820",
		16#2010# => X"d4016024",
		16#2011# => X"0400156d",
		16#2012# => X"a86385a9",
		16#2013# => X"18800001",
		16#2014# => X"84700008",
		16#2015# => X"84d00000",
		16#2016# => X"84b00004",
		16#2017# => X"a88485d7",
		16#2018# => X"87100010",
		16#2019# => X"d4013008",
		16#201a# => X"d401280c",
		16#201b# => X"d4011000",
		16#201c# => X"04000a6c",
		16#201d# => X"d4012004",
		16#201e# => X"8490000c",
		16#201f# => X"a8780000",
		16#2020# => X"d4015810",
		16#2021# => X"d4016014",
		16#2022# => X"d4012018",
		16#2023# => X"040009d8",
		16#2024# => X"d401c01c",
		16#2025# => X"18800001",
		16#2026# => X"84760000",
		16#2027# => X"a884bc48",
		16#2028# => X"ab0b0000",
		16#2029# => X"040009d2",
		16#202a# => X"e20e2000",
		16#202b# => X"18a00001",
		16#202c# => X"a88b0000",
		16#202d# => X"a8a5bcfc",
		16#202e# => X"a8780000",
		16#202f# => X"e0ae2800",
		16#2030# => X"04000820",
		16#2031# => X"d4012828",
		16#2032# => X"18c00001",
		16#2033# => X"a86b0000",
		16#2034# => X"a8c6bdb0",
		16#2035# => X"e0ce3000",
		16#2036# => X"04000a52",
		16#2037# => X"d4013034",
		16#2038# => X"18600001",
		16#2039# => X"d4015820",
		16#203a# => X"d4016024",
		16#203b# => X"04001543",
		16#203c# => X"a86385a9",
		16#203d# => X"18800001",
		16#203e# => X"84740008",
		16#203f# => X"84d40000",
		16#2040# => X"84b40004",
		16#2041# => X"a88485dd",
		16#2042# => X"87140010",
		16#2043# => X"d4013008",
		16#2044# => X"d401280c",
		16#2045# => X"d4011000",
		16#2046# => X"04000a42",
		16#2047# => X"d4012004",
		16#2048# => X"8494000c",
		16#2049# => X"a8780000",
		16#204a# => X"d4015810",
		16#204b# => X"d4016014",
		16#204c# => X"d4012018",
		16#204d# => X"040009ae",
		16#204e# => X"d401c01c",
		16#204f# => X"18800001",
		16#2050# => X"84760000",
		16#2051# => X"a884be64",
		16#2052# => X"ab0b0000",
		16#2053# => X"040009a8",
		16#2054# => X"e28e2000",
		16#2055# => X"18a00001",
		16#2056# => X"a88b0000",
		16#2057# => X"a8a5bf18",
		16#2058# => X"a8780000",
		16#2059# => X"e0ae2800",
		16#205a# => X"040007f6",
		16#205b# => X"d4012838",
		16#205c# => X"18c00001",
		16#205d# => X"a86b0000",
		16#205e# => X"a8c6bfcc",
		16#205f# => X"04000a29",
		16#2060# => X"e3ce3000",
		16#2061# => X"18600001",
		16#2062# => X"d4015820",
		16#2063# => X"d4016024",
		16#2064# => X"0400151a",
		16#2065# => X"a86385a9",
		16#2066# => X"18800001",
		16#2067# => X"84720008",
		16#2068# => X"84d20000",
		16#2069# => X"84b20004",
		16#206a# => X"a884874f",
		16#206b# => X"87120010",
		16#206c# => X"d4013008",
		16#206d# => X"d401280c",
		16#206e# => X"d4011000",
		16#206f# => X"04000a19",
		16#2070# => X"d4012004",
		16#2071# => X"8492000c",
		16#2072# => X"a8780000",
		16#2073# => X"d4015810",
		16#2074# => X"d4016014",
		16#2075# => X"d4012018",
		16#2076# => X"04000985",
		16#2077# => X"d401c01c",
		16#2078# => X"18800001",
		16#2079# => X"84760000",
		16#207a# => X"a884c080",
		16#207b# => X"ab0b0000",
		16#207c# => X"0400097f",
		16#207d# => X"e38e2000",
		16#207e# => X"18a00001",
		16#207f# => X"a88b0000",
		16#2080# => X"a8a5c134",
		16#2081# => X"a8780000",
		16#2082# => X"040007ce",
		16#2083# => X"e34e2800",
		16#2084# => X"18c00001",
		16#2085# => X"a86b0000",
		16#2086# => X"a8c6c1e8",
		16#2087# => X"04000a01",
		16#2088# => X"e30e3000",
		16#2089# => X"18600001",
		16#208a# => X"d4015820",
		16#208b# => X"d4016024",
		16#208c# => X"040014f2",
		16#208d# => X"a86385a9",
		16#208e# => X"18800001",
		16#208f# => X"84700008",
		16#2090# => X"84d00000",
		16#2091# => X"84b00004",
		16#2092# => X"a8848759",
		16#2093# => X"d4013008",
		16#2094# => X"d401280c",
		16#2095# => X"d4011000",
		16#2096# => X"040009f2",
		16#2097# => X"d4012004",
		16#2098# => X"8490000c",
		16#2099# => X"84700010",
		16#209a# => X"d4015810",
		16#209b# => X"d4016014",
		16#209c# => X"d4012018",
		16#209d# => X"0400095e",
		16#209e# => X"d401181c",
		16#209f# => X"18a00001",
		16#20a0# => X"84760000",
		16#20a1# => X"a8a5c29c",
		16#20a2# => X"d401582c",
		16#20a3# => X"04000958",
		16#20a4# => X"e1ce2800",
		16#20a5# => X"8461002c",
		16#20a6# => X"040007aa",
		16#20a7# => X"a88b0000",
		16#20a8# => X"040009e0",
		16#20a9# => X"a86b0000",
		16#20aa# => X"18600001",
		16#20ab# => X"d4015820",
		16#20ac# => X"d4016024",
		16#20ad# => X"040014d1",
		16#20ae# => X"a86385a9",
		16#20af# => X"84810028",
		16#20b0# => X"84c10028",
		16#20b1# => X"84a40004",
		16#20b2# => X"84840010",
		16#20b3# => X"84660008",
		16#20b4# => X"84c60000",
		16#20b5# => X"d401201c",
		16#20b6# => X"18800001",
		16#20b7# => X"d4013008",
		16#20b8# => X"a88485e1",
		16#20b9# => X"d4011000",
		16#20ba# => X"d4012004",
		16#20bb# => X"040009cd",
		16#20bc# => X"d401280c",
		16#20bd# => X"84a10028",
		16#20be# => X"8461001c",
		16#20bf# => X"8485000c",
		16#20c0# => X"d4015810",
		16#20c1# => X"d4016014",
		16#20c2# => X"04000939",
		16#20c3# => X"d4012018",
		16#20c4# => X"84760000",
		16#20c5# => X"04000936",
		16#20c6# => X"d4015828",
		16#20c7# => X"84610028",
		16#20c8# => X"04000788",
		16#20c9# => X"a88b0000",
		16#20ca# => X"040009be",
		16#20cb# => X"a86b0000",
		16#20cc# => X"18600001",
		16#20cd# => X"d4015820",
		16#20ce# => X"d4016024",
		16#20cf# => X"040014af",
		16#20d0# => X"a86385a9",
		16#20d1# => X"84810034",
		16#20d2# => X"84c10034",
		16#20d3# => X"84a40004",
		16#20d4# => X"84840010",
		16#20d5# => X"84660008",
		16#20d6# => X"84c60000",
		16#20d7# => X"d401201c",
		16#20d8# => X"18800001",
		16#20d9# => X"d4013008",
		16#20da# => X"a88485e6",
		16#20db# => X"d4011000",
		16#20dc# => X"d4012004",
		16#20dd# => X"040009ab",
		16#20de# => X"d401280c",
		16#20df# => X"84a10034",
		16#20e0# => X"8461001c",
		16#20e1# => X"8485000c",
		16#20e2# => X"d4015810",
		16#20e3# => X"d4016014",
		16#20e4# => X"04000917",
		16#20e5# => X"d4012018",
		16#20e6# => X"84760000",
		16#20e7# => X"04000914",
		16#20e8# => X"d4015828",
		16#20e9# => X"84610028",
		16#20ea# => X"04000766",
		16#20eb# => X"a88b0000",
		16#20ec# => X"0400099c",
		16#20ed# => X"a86b0000",
		16#20ee# => X"18600001",
		16#20ef# => X"d4015820",
		16#20f0# => X"d4016024",
		16#20f1# => X"0400148d",
		16#20f2# => X"a86385a9",
		16#20f3# => X"84810030",
		16#20f4# => X"84c10030",
		16#20f5# => X"84a40004",
		16#20f6# => X"18800001",
		16#20f7# => X"84660008",
		16#20f8# => X"a8848610",
		16#20f9# => X"84c60000",
		16#20fa# => X"d4011000",
		16#20fb# => X"d4012004",
		16#20fc# => X"d4013008",
		16#20fd# => X"0400098b",
		16#20fe# => X"d401280c",
		16#20ff# => X"84c10030",
		16#2100# => X"18600001",
		16#2101# => X"84a6000c",
		16#2102# => X"84960000",
		16#2103# => X"a86385ec",
		16#2104# => X"d4015810",
		16#2105# => X"d4016014",
		16#2106# => X"d4012818",
		16#2107# => X"04001477",
		16#2108# => X"d401201c",
		16#2109# => X"18800001",
		16#210a# => X"84740008",
		16#210b# => X"84d40000",
		16#210c# => X"84b40004",
		16#210d# => X"a8848617",
		16#210e# => X"d4013008",
		16#210f# => X"d4011000",
		16#2110# => X"d4012004",
		16#2111# => X"04000977",
		16#2112# => X"d401280c",
		16#2113# => X"18600001",
		16#2114# => X"84b4000c",
		16#2115# => X"84940010",
		16#2116# => X"a86385ec",
		16#2117# => X"d4015810",
		16#2118# => X"d4016014",
		16#2119# => X"d4012818",
		16#211a# => X"04001464",
		16#211b# => X"d401201c",
		16#211c# => X"84810038",
		16#211d# => X"84640008",
		16#211e# => X"86c40000",
		16#211f# => X"84a40004",
		16#2120# => X"18800001",
		16#2121# => X"d4011000",
		16#2122# => X"a8848614",
		16#2123# => X"d401b008",
		16#2124# => X"d4012004",
		16#2125# => X"04000963",
		16#2126# => X"d401280c",
		16#2127# => X"84c10038",
		16#2128# => X"a8760000",
		16#2129# => X"84a6000c",
		16#212a# => X"84860010",
		16#212b# => X"d4012818",
		16#212c# => X"d4015810",
		16#212d# => X"d4016014",
		16#212e# => X"040008cd",
		16#212f# => X"d401201c",
		16#2130# => X"84740000",
		16#2131# => X"040008ca",
		16#2132# => X"aacb0000",
		16#2133# => X"a8760000",
		16#2134# => X"0400071c",
		16#2135# => X"a88b0000",
		16#2136# => X"04000952",
		16#2137# => X"a86b0000",
		16#2138# => X"18600001",
		16#2139# => X"d4015820",
		16#213a# => X"d4016024",
		16#213b# => X"04001443",
		16#213c# => X"a86385a9",
		16#213d# => X"18800001",
		16#213e# => X"847e0008",
		16#213f# => X"86de0000",
		16#2140# => X"84be0004",
		16#2141# => X"a884861b",
		16#2142# => X"d4011000",
		16#2143# => X"d4012004",
		16#2144# => X"d401b008",
		16#2145# => X"04000943",
		16#2146# => X"d401280c",
		16#2147# => X"84be000c",
		16#2148# => X"849e0010",
		16#2149# => X"a8760000",
		16#214a# => X"d4012818",
		16#214b# => X"d4015810",
		16#214c# => X"d4016014",
		16#214d# => X"040008ae",
		16#214e# => X"d401201c",
		16#214f# => X"84740000",
		16#2150# => X"040008ab",
		16#2151# => X"aacb0000",
		16#2152# => X"a8760000",
		16#2153# => X"040006fd",
		16#2154# => X"a88b0000",
		16#2155# => X"04000933",
		16#2156# => X"a86b0000",
		16#2157# => X"18600001",
		16#2158# => X"d4015820",
		16#2159# => X"d4016024",
		16#215a# => X"04001424",
		16#215b# => X"a86385a9",
		16#215c# => X"18800001",
		16#215d# => X"847c0008",
		16#215e# => X"869c0000",
		16#215f# => X"84bc0004",
		16#2160# => X"a8848622",
		16#2161# => X"d4011000",
		16#2162# => X"d4012004",
		16#2163# => X"d401a008",
		16#2164# => X"04000924",
		16#2165# => X"d401280c",
		16#2166# => X"84bc000c",
		16#2167# => X"849c0010",
		16#2168# => X"a8740000",
		16#2169# => X"d4012818",
		16#216a# => X"d4015810",
		16#216b# => X"d4016014",
		16#216c# => X"0400088f",
		16#216d# => X"d401201c",
		16#216e# => X"84720000",
		16#216f# => X"0400088c",
		16#2170# => X"aa8b0000",
		16#2171# => X"a8740000",
		16#2172# => X"040006de",
		16#2173# => X"a88b0000",
		16#2174# => X"04000914",
		16#2175# => X"a86b0000",
		16#2176# => X"18600001",
		16#2177# => X"d4015820",
		16#2178# => X"d4016024",
		16#2179# => X"04001405",
		16#217a# => X"a86385a9",
		16#217b# => X"18800001",
		16#217c# => X"847a0008",
		16#217d# => X"869a0000",
		16#217e# => X"84ba0004",
		16#217f# => X"a8848629",
		16#2180# => X"d4011000",
		16#2181# => X"d4012004",
		16#2182# => X"d401a008",
		16#2183# => X"04000905",
		16#2184# => X"d401280c",
		16#2185# => X"84ba000c",
		16#2186# => X"849a0010",
		16#2187# => X"a8740000",
		16#2188# => X"d4012818",
		16#2189# => X"d4015810",
		16#218a# => X"d4016014",
		16#218b# => X"04000870",
		16#218c# => X"d401201c",
		16#218d# => X"84720000",
		16#218e# => X"0400086d",
		16#218f# => X"aa8b0000",
		16#2190# => X"a8740000",
		16#2191# => X"040006bf",
		16#2192# => X"a88b0000",
		16#2193# => X"040008f5",
		16#2194# => X"a86b0000",
		16#2195# => X"18600001",
		16#2196# => X"d4015820",
		16#2197# => X"d4016024",
		16#2198# => X"040013e6",
		16#2199# => X"a86385a9",
		16#219a# => X"18800001",
		16#219b# => X"84780008",
		16#219c# => X"86580000",
		16#219d# => X"84b80004",
		16#219e# => X"a8848630",
		16#219f# => X"d4011000",
		16#21a0# => X"d4012004",
		16#21a1# => X"d4019008",
		16#21a2# => X"040008e6",
		16#21a3# => X"d401280c",
		16#21a4# => X"84b8000c",
		16#21a5# => X"84980010",
		16#21a6# => X"a8720000",
		16#21a7# => X"d4012818",
		16#21a8# => X"d4015810",
		16#21a9# => X"d4016014",
		16#21aa# => X"04000851",
		16#21ab# => X"d401201c",
		16#21ac# => X"84700000",
		16#21ad# => X"0400084e",
		16#21ae# => X"aa4b0000",
		16#21af# => X"a8720000",
		16#21b0# => X"040006a0",
		16#21b1# => X"a88b0000",
		16#21b2# => X"040008d6",
		16#21b3# => X"a86b0000",
		16#21b4# => X"18600001",
		16#21b5# => X"d4015820",
		16#21b6# => X"d4016024",
		16#21b7# => X"040013c7",
		16#21b8# => X"a86385a9",
		16#21b9# => X"846e0008",
		16#21ba# => X"864e0000",
		16#21bb# => X"848e0004",
		16#21bc# => X"d4011000",
		16#21bd# => X"18400001",
		16#21be# => X"d4019008",
		16#21bf# => X"a8428637",
		16#21c0# => X"d401200c",
		16#21c1# => X"040008c7",
		16#21c2# => X"d4011004",
		16#21c3# => X"848e000c",
		16#21c4# => X"844e0010",
		16#21c5# => X"a8720000",
		16#21c6# => X"d4015810",
		16#21c7# => X"d4016014",
		16#21c8# => X"d4012018",
		16#21c9# => X"04000832",
		16#21ca# => X"d401101c",
		16#21cb# => X"84700000",
		16#21cc# => X"0400082f",
		16#21cd# => X"a84b0000",
		16#21ce# => X"a8620000",
		16#21cf# => X"04000681",
		16#21d0# => X"a88b0000",
		16#21d1# => X"040008b7",
		16#21d2# => X"a86b0000",
		16#21d3# => X"18600001",
		16#21d4# => X"d4015820",
		16#21d5# => X"d4016024",
		16#21d6# => X"040013a8",
		16#21d7# => X"a86385a9",
		16#21d8# => X"9c210068",
		16#21d9# => X"8521fffc",
		16#21da# => X"8441ffd4",
		16#21db# => X"85c1ffd8",
		16#21dc# => X"8601ffdc",
		16#21dd# => X"8641ffe0",
		16#21de# => X"8681ffe4",
		16#21df# => X"86c1ffe8",
		16#21e0# => X"8701ffec",
		16#21e1# => X"8741fff0",
		16#21e2# => X"8781fff4",
		16#21e3# => X"44004800",
		16#21e4# => X"87c1fff8",
		16#21e5# => X"d7e177f8",
		16#21e6# => X"d7e14ffc",
		16#21e7# => X"d7e117f4",
		16#21e8# => X"9c21fff4",
		16#21e9# => X"040003aa",
		16#21ea# => X"a9c30000",
		16#21eb# => X"bc0b0000",
		16#21ec# => X"10000031",
		16#21ed# => X"9ca00000",
		16#21ee# => X"18c00fff",
		16#21ef# => X"9c8e0004",
		16#21f0# => X"a8c6ffff",
		16#21f1# => X"a8450000",
		16#21f2# => X"84e40000",
		16#21f3# => X"e4a63800",
		16#21f4# => X"10000003",
		16#21f5# => X"9c420001",
		16#21f6# => X"a8c70000",
		16#21f7# => X"84e40008",
		16#21f8# => X"e4653800",
		16#21f9# => X"10000003",
		16#21fa# => X"9c840014",
		16#21fb# => X"a8a70000",
		16#21fc# => X"e4825800",
		16#21fd# => X"13fffff5",
		16#21fe# => X"a86e0000",
		16#21ff# => X"9c4e00a0",
		16#2200# => X"d4023004",
		16#2201# => X"d402280c",
		16#2202# => X"84c20010",
		16#2203# => X"84a20000",
		16#2204# => X"9c800000",
		16#2205# => X"85030010",
		16#2206# => X"84e30000",
		16#2207# => X"e0c64000",
		16#2208# => X"e0a53800",
		16#2209# => X"9c840001",
		16#220a# => X"d4023010",
		16#220b# => X"d4022800",
		16#220c# => X"e44b2000",
		16#220d# => X"13fffff8",
		16#220e# => X"9c630014",
		16#220f# => X"040007ec",
		16#2210# => X"84620010",
		16#2211# => X"84620000",
		16#2212# => X"040007e9",
		16#2213# => X"a9cb0000",
		16#2214# => X"a86e0000",
		16#2215# => X"0400063b",
		16#2216# => X"a88b0000",
		16#2217# => X"d4025808",
		16#2218# => X"9c21000c",
		16#2219# => X"8521fffc",
		16#221a# => X"8441fff4",
		16#221b# => X"44004800",
		16#221c# => X"85c1fff8",
		16#221d# => X"18600fff",
		16#221e# => X"9c4e00a0",
		16#221f# => X"a863ffff",
		16#2220# => X"d402580c",
		16#2221# => X"03ffffee",
		16#2222# => X"d4021804",
		16#2223# => X"18600001",
		16#2224# => X"d7e14ffc",
		16#2225# => X"d7e117f0",
		16#2226# => X"d7e177f4",
		16#2227# => X"d7e187f8",
		16#2228# => X"a863b8c4",
		16#2229# => X"9c21fff0",
		16#222a# => X"07ffffbb",
		16#222b# => X"18400001",
		16#222c# => X"18600001",
		16#222d# => X"a842b978",
		16#222e# => X"07ffffb7",
		16#222f# => X"a863ba2c",
		16#2230# => X"18600001",
		16#2231# => X"07ffffb4",
		16#2232# => X"a863bae0",
		16#2233# => X"18600001",
		16#2234# => X"07ffffb1",
		16#2235# => X"a863bb94",
		16#2236# => X"18600001",
		16#2237# => X"07ffffae",
		16#2238# => X"a863bc48",
		16#2239# => X"18600001",
		16#223a# => X"07ffffab",
		16#223b# => X"a863bcfc",
		16#223c# => X"18600001",
		16#223d# => X"07ffffa8",
		16#223e# => X"a863bdb0",
		16#223f# => X"18600001",
		16#2240# => X"07ffffa5",
		16#2241# => X"a863be64",
		16#2242# => X"18600001",
		16#2243# => X"07ffffa2",
		16#2244# => X"a863c350",
		16#2245# => X"18600001",
		16#2246# => X"07ffff9f",
		16#2247# => X"a863c404",
		16#2248# => X"18600001",
		16#2249# => X"07ffff9c",
		16#224a# => X"a863bf18",
		16#224b# => X"18600001",
		16#224c# => X"07ffff99",
		16#224d# => X"a863bfcc",
		16#224e# => X"18600001",
		16#224f# => X"07ffff96",
		16#2250# => X"a863c080",
		16#2251# => X"18600001",
		16#2252# => X"07ffff93",
		16#2253# => X"a863c134",
		16#2254# => X"18600001",
		16#2255# => X"07ffff90",
		16#2256# => X"a863c1e8",
		16#2257# => X"18600001",
		16#2258# => X"07ffff8d",
		16#2259# => X"a863c29c",
		16#225a# => X"18c00001",
		16#225b# => X"18800001",
		16#225c# => X"a8c6ba2c",
		16#225d# => X"a884b8c4",
		16#225e# => X"18a00001",
		16#225f# => X"846400b0",
		16#2260# => X"84e600b0",
		16#2261# => X"a8a5bae0",
		16#2262# => X"e0e71800",
		16#2263# => X"850500b0",
		16#2264# => X"85c600a0",
		16#2265# => X"18600001",
		16#2266# => X"84c400a0",
		16#2267# => X"84a500a0",
		16#2268# => X"e0874000",
		16#2269# => X"a863bb94",
		16#226a# => X"e1ce3000",
		16#226b# => X"18e00001",
		16#226c# => X"850300b0",
		16#226d# => X"a8e7bc48",
		16#226e# => X"846300a0",
		16#226f# => X"e1ce2800",
		16#2270# => X"18c00001",
		16#2271# => X"e0844000",
		16#2272# => X"a8c6bcfc",
		16#2273# => X"850700b0",
		16#2274# => X"e1ce1800",
		16#2275# => X"18a00001",
		16#2276# => X"846700a0",
		16#2277# => X"e0844000",
		16#2278# => X"a8a5bdb0",
		16#2279# => X"850600b0",
		16#227a# => X"e1ce1800",
		16#227b# => X"846600a0",
		16#227c# => X"84e500b0",
		16#227d# => X"e0844000",
		16#227e# => X"84a500a0",
		16#227f# => X"e1ce1800",
		16#2280# => X"e0843800",
		16#2281# => X"e1ce2800",
		16#2282# => X"a8640000",
		16#2283# => X"d40220b0",
		16#2284# => X"04000777",
		16#2285# => X"d40270a0",
		16#2286# => X"a86e0000",
		16#2287# => X"04000774",
		16#2288# => X"aa0b0000",
		16#2289# => X"a8700000",
		16#228a# => X"040005c6",
		16#228b# => X"a88b0000",
		16#228c# => X"d40258a8",
		16#228d# => X"9c210010",
		16#228e# => X"8521fffc",
		16#228f# => X"8441fff0",
		16#2290# => X"85c1fff4",
		16#2291# => X"44004800",
		16#2292# => X"8601fff8",
		16#2293# => X"18600001",
		16#2294# => X"d7e14ffc",
		16#2295# => X"d7e117d4",
		16#2296# => X"d7e177d8",
		16#2297# => X"d7e187dc",
		16#2298# => X"d7e197e0",
		16#2299# => X"d7e1a7e4",
		16#229a# => X"d7e1b7e8",
		16#229b# => X"d7e1c7ec",
		16#229c# => X"d7e1d7f0",
		16#229d# => X"d7e1e7f4",
		16#229e# => X"d7e1f7f8",
		16#229f# => X"a863863e",
		16#22a0# => X"9c21ffac",
		16#22a1# => X"040013c0",
		16#22a2# => X"19c00001",
		16#22a3# => X"18600001",
		16#22a4# => X"a9ceb8c4",
		16#22a5# => X"a8638688",
		16#22a6# => X"040013bb",
		16#22a7# => X"18400001",
		16#22a8# => X"18800001",
		16#22a9# => X"18600001",
		16#22aa# => X"a8848586",
		16#22ab# => X"a86386b1",
		16#22ac# => X"d4012000",
		16#22ad# => X"18800001",
		16#22ae# => X"a842b978",
		16#22af# => X"a884858c",
		16#22b0# => X"1a400001",
		16#22b1# => X"d4012004",
		16#22b2# => X"18800001",
		16#22b3# => X"aa52ba2c",
		16#22b4# => X"a8848592",
		16#22b5# => X"1a800001",
		16#22b6# => X"d4012008",
		16#22b7# => X"18800001",
		16#22b8# => X"aa94bae0",
		16#22b9# => X"a8848596",
		16#22ba# => X"1bc00001",
		16#22bb# => X"d401200c",
		16#22bc# => X"18800001",
		16#22bd# => X"abdec080",
		16#22be# => X"a884859a",
		16#22bf# => X"1b800001",
		16#22c0# => X"d4012010",
		16#22c1# => X"18800001",
		16#22c2# => X"ab9cc134",
		16#22c3# => X"a884859e",
		16#22c4# => X"1b400001",
		16#22c5# => X"d4012014",
		16#22c6# => X"18800001",
		16#22c7# => X"ab5ac1e8",
		16#22c8# => X"a88485a4",
		16#22c9# => X"1b000001",
		16#22ca# => X"040012b4",
		16#22cb# => X"d4012018",
		16#22cc# => X"18600001",
		16#22cd# => X"ab18c29c",
		16#22ce# => X"04001393",
		16#22cf# => X"a863863e",
		16#22d0# => X"18800001",
		16#22d1# => X"846e00a8",
		16#22d2# => X"84ce00a0",
		16#22d3# => X"84ae00a4",
		16#22d4# => X"a88485d3",
		16#22d5# => X"860e00b0",
		16#22d6# => X"d4013004",
		16#22d7# => X"d4012808",
		16#22d8# => X"040007b0",
		16#22d9# => X"d4012000",
		16#22da# => X"848e00ac",
		16#22db# => X"a8700000",
		16#22dc# => X"d401580c",
		16#22dd# => X"d4016010",
		16#22de# => X"d4012014",
		16#22df# => X"0400071c",
		16#22e0# => X"d4018018",
		16#22e1# => X"846200b0",
		16#22e2# => X"04000719",
		16#22e3# => X"a9cb0000",
		16#22e4# => X"a86e0000",
		16#22e5# => X"a88b0000",
		16#22e6# => X"0400056a",
		16#22e7# => X"1a000001",
		16#22e8# => X"a86b0000",
		16#22e9# => X"0400079f",
		16#22ea# => X"aa10bb94",
		16#22eb# => X"18600001",
		16#22ec# => X"d401581c",
		16#22ed# => X"d4016020",
		16#22ee# => X"a86386d6",
		16#22ef# => X"0400128f",
		16#22f0# => X"19c00001",
		16#22f1# => X"18800001",
		16#22f2# => X"847200a8",
		16#22f3# => X"84d200a0",
		16#22f4# => X"84b200a4",
		16#22f5# => X"a88485d7",
		16#22f6# => X"86d200b0",
		16#22f7# => X"d4013004",
		16#22f8# => X"d4012808",
		16#22f9# => X"0400078f",
		16#22fa# => X"d4012000",
		16#22fb# => X"849200ac",
		16#22fc# => X"a8760000",
		16#22fd# => X"d401580c",
		16#22fe# => X"d4016010",
		16#22ff# => X"d4012014",
		16#2300# => X"040006fb",
		16#2301# => X"d401b018",
		16#2302# => X"846200b0",
		16#2303# => X"040006f8",
		16#2304# => X"aa4b0000",
		16#2305# => X"a8720000",
		16#2306# => X"a88b0000",
		16#2307# => X"04000549",
		16#2308# => X"a9cebc48",
		16#2309# => X"a86b0000",
		16#230a# => X"0400077e",
		16#230b# => X"1a400001",
		16#230c# => X"18600001",
		16#230d# => X"d401581c",
		16#230e# => X"d4016020",
		16#230f# => X"a86386d6",
		16#2310# => X"0400126e",
		16#2311# => X"aa52be64",
		16#2312# => X"18800001",
		16#2313# => X"847400a8",
		16#2314# => X"84d400a0",
		16#2315# => X"84b400a4",
		16#2316# => X"a88485dd",
		16#2317# => X"86d400b0",
		16#2318# => X"d4013004",
		16#2319# => X"d4012808",
		16#231a# => X"0400076e",
		16#231b# => X"d4012000",
		16#231c# => X"849400ac",
		16#231d# => X"a8760000",
		16#231e# => X"d401580c",
		16#231f# => X"d4016010",
		16#2320# => X"d4012014",
		16#2321# => X"040006da",
		16#2322# => X"d401b018",
		16#2323# => X"846200b0",
		16#2324# => X"040006d7",
		16#2325# => X"aa8b0000",
		16#2326# => X"a8740000",
		16#2327# => X"a88b0000",
		16#2328# => X"04000528",
		16#2329# => X"1ac00001",
		16#232a# => X"a86b0000",
		16#232b# => X"0400075d",
		16#232c# => X"aad6c350",
		16#232d# => X"18600001",
		16#232e# => X"d401581c",
		16#232f# => X"d4016020",
		16#2330# => X"0400124e",
		16#2331# => X"a86386d6",
		16#2332# => X"18800001",
		16#2333# => X"847000a8",
		16#2334# => X"84d000a0",
		16#2335# => X"84b000a4",
		16#2336# => X"a884874f",
		16#2337# => X"869000b0",
		16#2338# => X"d4013004",
		16#2339# => X"d4012808",
		16#233a# => X"0400074e",
		16#233b# => X"d4012000",
		16#233c# => X"849000ac",
		16#233d# => X"a8740000",
		16#233e# => X"d401580c",
		16#233f# => X"d4016010",
		16#2340# => X"d4012014",
		16#2341# => X"040006ba",
		16#2342# => X"d401a018",
		16#2343# => X"846200b0",
		16#2344# => X"040006b7",
		16#2345# => X"aa8b0000",
		16#2346# => X"a8740000",
		16#2347# => X"04000509",
		16#2348# => X"a88b0000",
		16#2349# => X"0400073f",
		16#234a# => X"a86b0000",
		16#234b# => X"18600001",
		16#234c# => X"d401581c",
		16#234d# => X"d4016020",
		16#234e# => X"04001230",
		16#234f# => X"a86386d6",
		16#2350# => X"18800001",
		16#2351# => X"846e00a8",
		16#2352# => X"84ce00a0",
		16#2353# => X"84ae00a4",
		16#2354# => X"a8848759",
		16#2355# => X"868e00b0",
		16#2356# => X"d4013004",
		16#2357# => X"d4012808",
		16#2358# => X"04000730",
		16#2359# => X"d4012000",
		16#235a# => X"848e00ac",
		16#235b# => X"a8740000",
		16#235c# => X"d401580c",
		16#235d# => X"d4016010",
		16#235e# => X"d4012014",
		16#235f# => X"0400069c",
		16#2360# => X"d401a018",
		16#2361# => X"846200b0",
		16#2362# => X"04000699",
		16#2363# => X"aa8b0000",
		16#2364# => X"a8740000",
		16#2365# => X"a88b0000",
		16#2366# => X"040004ea",
		16#2367# => X"1a800001",
		16#2368# => X"a86b0000",
		16#2369# => X"0400071f",
		16#236a# => X"aa94c404",
		16#236b# => X"18600001",
		16#236c# => X"d401581c",
		16#236d# => X"d4016020",
		16#236e# => X"04001210",
		16#236f# => X"a86386d6",
		16#2370# => X"18800001",
		16#2371# => X"a884bcfc",
		16#2372# => X"84c400a0",
		16#2373# => X"846400a8",
		16#2374# => X"84a400a4",
		16#2375# => X"848400b0",
		16#2376# => X"d4013004",
		16#2377# => X"d4012018",
		16#2378# => X"18800001",
		16#2379# => X"d4012808",
		16#237a# => X"a88485e1",
		16#237b# => X"0400070d",
		16#237c# => X"d4012000",
		16#237d# => X"18a00001",
		16#237e# => X"84610018",
		16#237f# => X"a8a5bcfc",
		16#2380# => X"848500ac",
		16#2381# => X"d401580c",
		16#2382# => X"d4016010",
		16#2383# => X"04000678",
		16#2384# => X"d4012014",
		16#2385# => X"846200b0",
		16#2386# => X"04000675",
		16#2387# => X"d4015824",
		16#2388# => X"84610024",
		16#2389# => X"040004c7",
		16#238a# => X"a88b0000",
		16#238b# => X"040006fd",
		16#238c# => X"a86b0000",
		16#238d# => X"18600001",
		16#238e# => X"d401581c",
		16#238f# => X"d4016020",
		16#2390# => X"040011ee",
		16#2391# => X"a86386d6",
		16#2392# => X"18800001",
		16#2393# => X"a884bdb0",
		16#2394# => X"84c400a0",
		16#2395# => X"846400a8",
		16#2396# => X"84a400a4",
		16#2397# => X"848400b0",
		16#2398# => X"d4013004",
		16#2399# => X"d4012018",
		16#239a# => X"18800001",
		16#239b# => X"d4012808",
		16#239c# => X"a88485e6",
		16#239d# => X"040006eb",
		16#239e# => X"d4012000",
		16#239f# => X"18a00001",
		16#23a0# => X"84610018",
		16#23a1# => X"a8a5bdb0",
		16#23a2# => X"848500ac",
		16#23a3# => X"d401580c",
		16#23a4# => X"d4016010",
		16#23a5# => X"04000656",
		16#23a6# => X"d4012014",
		16#23a7# => X"846200b0",
		16#23a8# => X"04000653",
		16#23a9# => X"d4015824",
		16#23aa# => X"84610024",
		16#23ab# => X"040004a5",
		16#23ac# => X"a88b0000",
		16#23ad# => X"040006db",
		16#23ae# => X"a86b0000",
		16#23af# => X"18600001",
		16#23b0# => X"d401581c",
		16#23b1# => X"d4016020",
		16#23b2# => X"040011cc",
		16#23b3# => X"a86386d6",
		16#23b4# => X"848200a0",
		16#23b5# => X"84a200a4",
		16#23b6# => X"846200a8",
		16#23b7# => X"d4012004",
		16#23b8# => X"18800001",
		16#23b9# => X"d4012808",
		16#23ba# => X"a8848610",
		16#23bb# => X"040006cd",
		16#23bc# => X"d4012000",
		16#23bd# => X"18600001",
		16#23be# => X"848200ac",
		16#23bf# => X"a86386ff",
		16#23c0# => X"844200b0",
		16#23c1# => X"d401580c",
		16#23c2# => X"d4016010",
		16#23c3# => X"d4012014",
		16#23c4# => X"040011ba",
		16#23c5# => X"d4011018",
		16#23c6# => X"845200a0",
		16#23c7# => X"847200a8",
		16#23c8# => X"849200a4",
		16#23c9# => X"d4011004",
		16#23ca# => X"18400001",
		16#23cb# => X"d4012008",
		16#23cc# => X"a8428617",
		16#23cd# => X"040006bb",
		16#23ce# => X"d4011000",
		16#23cf# => X"18600001",
		16#23d0# => X"849200ac",
		16#23d1# => X"845200b0",
		16#23d2# => X"a86386ff",
		16#23d3# => X"d401580c",
		16#23d4# => X"d4016010",
		16#23d5# => X"d4012014",
		16#23d6# => X"040011a8",
		16#23d7# => X"d4011018",
		16#23d8# => X"18800001",
		16#23d9# => X"18400001",
		16#23da# => X"a884bf18",
		16#23db# => X"a842bf18",
		16#23dc# => X"84a400a4",
		16#23dd# => X"18800001",
		16#23de# => X"846200a8",
		16#23df# => X"a8848614",
		16#23e0# => X"844200a0",
		16#23e1# => X"d4012000",
		16#23e2# => X"d4011004",
		16#23e3# => X"040006a5",
		16#23e4# => X"d4012808",
		16#23e5# => X"18a00001",
		16#23e6# => X"a8620000",
		16#23e7# => X"a8a5bf18",
		16#23e8# => X"848500ac",
		16#23e9# => X"844500b0",
		16#23ea# => X"d401580c",
		16#23eb# => X"d4016010",
		16#23ec# => X"d4012014",
		16#23ed# => X"0400060e",
		16#23ee# => X"d4011018",
		16#23ef# => X"847200a0",
		16#23f0# => X"0400060b",
		16#23f1# => X"a84b0000",
		16#23f2# => X"a8620000",
		16#23f3# => X"a88b0000",
		16#23f4# => X"0400045c",
		16#23f5# => X"18400001",
		16#23f6# => X"a86b0000",
		16#23f7# => X"04000691",
		16#23f8# => X"a842bfcc",
		16#23f9# => X"18600001",
		16#23fa# => X"d401581c",
		16#23fb# => X"d4016020",
		16#23fc# => X"04001182",
		16#23fd# => X"a86386d6",
		16#23fe# => X"18800001",
		16#23ff# => X"846200a8",
		16#2400# => X"a884bfcc",
		16#2401# => X"844200a0",
		16#2402# => X"84a400a4",
		16#2403# => X"18800001",
		16#2404# => X"d4011004",
		16#2405# => X"a884861b",
		16#2406# => X"d4012808",
		16#2407# => X"04000681",
		16#2408# => X"d4012000",
		16#2409# => X"18a00001",
		16#240a# => X"a8620000",
		16#240b# => X"a8a5bfcc",
		16#240c# => X"848500ac",
		16#240d# => X"844500b0",
		16#240e# => X"d401580c",
		16#240f# => X"d4016010",
		16#2410# => X"d4012014",
		16#2411# => X"040005ea",
		16#2412# => X"d4011018",
		16#2413# => X"847200a0",
		16#2414# => X"040005e7",
		16#2415# => X"a84b0000",
		16#2416# => X"a8620000",
		16#2417# => X"04000439",
		16#2418# => X"a88b0000",
		16#2419# => X"0400066f",
		16#241a# => X"a86b0000",
		16#241b# => X"18600001",
		16#241c# => X"d401581c",
		16#241d# => X"d4016020",
		16#241e# => X"04001160",
		16#241f# => X"a86386d6",
		16#2420# => X"18800001",
		16#2421# => X"847e00a8",
		16#2422# => X"84be00a4",
		16#2423# => X"845e00a0",
		16#2424# => X"a8848622",
		16#2425# => X"d4012808",
		16#2426# => X"d4011004",
		16#2427# => X"04000661",
		16#2428# => X"d4012000",
		16#2429# => X"849e00ac",
		16#242a# => X"a8620000",
		16#242b# => X"845e00b0",
		16#242c# => X"d401580c",
		16#242d# => X"d4016010",
		16#242e# => X"d4012014",
		16#242f# => X"040005cc",
		16#2430# => X"d4011018",
		16#2431# => X"847000a0",
		16#2432# => X"040005c9",
		16#2433# => X"a84b0000",
		16#2434# => X"a8620000",
		16#2435# => X"0400041b",
		16#2436# => X"a88b0000",
		16#2437# => X"04000651",
		16#2438# => X"a86b0000",
		16#2439# => X"18600001",
		16#243a# => X"d401581c",
		16#243b# => X"d4016020",
		16#243c# => X"04001142",
		16#243d# => X"a86386d6",
		16#243e# => X"18800001",
		16#243f# => X"847c00a8",
		16#2440# => X"84bc00a4",
		16#2441# => X"845c00a0",
		16#2442# => X"a8848629",
		16#2443# => X"d4012808",
		16#2444# => X"d4011004",
		16#2445# => X"04000643",
		16#2446# => X"d4012000",
		16#2447# => X"849c00ac",
		16#2448# => X"a8620000",
		16#2449# => X"845c00b0",
		16#244a# => X"d401580c",
		16#244b# => X"d4016010",
		16#244c# => X"d4012014",
		16#244d# => X"040005ae",
		16#244e# => X"d4011018",
		16#244f# => X"847000a0",
		16#2450# => X"040005ab",
		16#2451# => X"a84b0000",
		16#2452# => X"a8620000",
		16#2453# => X"040003fd",
		16#2454# => X"a88b0000",
		16#2455# => X"04000633",
		16#2456# => X"a86b0000",
		16#2457# => X"18600001",
		16#2458# => X"d401581c",
		16#2459# => X"d4016020",
		16#245a# => X"04001124",
		16#245b# => X"a86386d6",
		16#245c# => X"18800001",
		16#245d# => X"847a00a8",
		16#245e# => X"84ba00a4",
		16#245f# => X"845a00a0",
		16#2460# => X"a8848630",
		16#2461# => X"d4012808",
		16#2462# => X"d4011004",
		16#2463# => X"04000625",
		16#2464# => X"d4012000",
		16#2465# => X"849a00ac",
		16#2466# => X"a8620000",
		16#2467# => X"845a00b0",
		16#2468# => X"d401580c",
		16#2469# => X"d4016010",
		16#246a# => X"d4012014",
		16#246b# => X"04000590",
		16#246c# => X"d4011018",
		16#246d# => X"846e00a0",
		16#246e# => X"0400058d",
		16#246f# => X"a84b0000",
		16#2470# => X"a8620000",
		16#2471# => X"040003df",
		16#2472# => X"a88b0000",
		16#2473# => X"04000615",
		16#2474# => X"a86b0000",
		16#2475# => X"18600001",
		16#2476# => X"d401581c",
		16#2477# => X"d4016020",
		16#2478# => X"04001106",
		16#2479# => X"a86386d6",
		16#247a# => X"18800001",
		16#247b# => X"847800a8",
		16#247c# => X"84b800a4",
		16#247d# => X"845800a0",
		16#247e# => X"a8848637",
		16#247f# => X"d4012808",
		16#2480# => X"d4011004",
		16#2481# => X"04000607",
		16#2482# => X"d4012000",
		16#2483# => X"849800ac",
		16#2484# => X"a8620000",
		16#2485# => X"845800b0",
		16#2486# => X"d401580c",
		16#2487# => X"d4016010",
		16#2488# => X"d4012014",
		16#2489# => X"04000572",
		16#248a# => X"d4011018",
		16#248b# => X"846e00a0",
		16#248c# => X"0400056f",
		16#248d# => X"a84b0000",
		16#248e# => X"a8620000",
		16#248f# => X"040003c1",
		16#2490# => X"a88b0000",
		16#2491# => X"040005f7",
		16#2492# => X"a86b0000",
		16#2493# => X"18600001",
		16#2494# => X"d401581c",
		16#2495# => X"d4016020",
		16#2496# => X"040010e8",
		16#2497# => X"a86386d6",
		16#2498# => X"84560000",
		16#2499# => X"84760008",
		16#249a# => X"84960004",
		16#249b# => X"d4011004",
		16#249c# => X"18400001",
		16#249d# => X"d4012008",
		16#249e# => X"a8428722",
		16#249f# => X"040005e9",
		16#24a0# => X"d4011000",
		16#24a1# => X"18600001",
		16#24a2# => X"8496000c",
		16#24a3# => X"84560010",
		16#24a4# => X"a86386ff",
		16#24a5# => X"d401580c",
		16#24a6# => X"d4016010",
		16#24a7# => X"d4012014",
		16#24a8# => X"040010d6",
		16#24a9# => X"d4011018",
		16#24aa# => X"18400001",
		16#24ab# => X"84740008",
		16#24ac# => X"84940004",
		16#24ad# => X"84b40000",
		16#24ae# => X"a8428726",
		16#24af# => X"d4012804",
		16#24b0# => X"d4011000",
		16#24b1# => X"040005d7",
		16#24b2# => X"d4012008",
		16#24b3# => X"18600001",
		16#24b4# => X"84540010",
		16#24b5# => X"8494000c",
		16#24b6# => X"a86386ff",
		16#24b7# => X"d4011018",
		16#24b8# => X"d401580c",
		16#24b9# => X"d4016010",
		16#24ba# => X"040010c4",
		16#24bb# => X"d4012014",
		16#24bc# => X"9c210054",
		16#24bd# => X"8521fffc",
		16#24be# => X"8441ffd4",
		16#24bf# => X"85c1ffd8",
		16#24c0# => X"8601ffdc",
		16#24c1# => X"8641ffe0",
		16#24c2# => X"8681ffe4",
		16#24c3# => X"86c1ffe8",
		16#24c4# => X"8701ffec",
		16#24c5# => X"8741fff0",
		16#24c6# => X"8781fff4",
		16#24c7# => X"44004800",
		16#24c8# => X"87c1fff8",
		16#24c9# => X"d7e177ec",
		16#24ca# => X"d7e187f0",
		16#24cb# => X"d7e197f4",
		16#24cc# => X"d7e14ffc",
		16#24cd# => X"d7e117e8",
		16#24ce# => X"d7e1a7f8",
		16#24cf# => X"a9c40000",
		16#24d0# => X"9c21ffd8",
		16#24d1# => X"aa030000",
		16#24d2# => X"bda40000",
		16#24d3# => X"10000012",
		16#24d4# => X"aa460000",
		16#24d5# => X"a860c7ff",
		16#24d6# => X"9c400000",
		16#24d7# => X"e2851800",
		16#24d8# => X"9c420001",
		16#24d9# => X"04001042",
		16#24da# => X"e0741000",
		16#24db# => X"18600001",
		16#24dc# => X"d4018000",
		16#24dd# => X"a863872b",
		16#24de# => X"d4019004",
		16#24df# => X"d4011008",
		16#24e0# => X"0400109e",
		16#24e1# => X"d401580c",
		16#24e2# => X"e54e1000",
		16#24e3# => X"13fffff6",
		16#24e4# => X"9c420001",
		16#24e5# => X"9c210028",
		16#24e6# => X"8521fffc",
		16#24e7# => X"8441ffe8",
		16#24e8# => X"85c1ffec",
		16#24e9# => X"8601fff0",
		16#24ea# => X"8641fff4",
		16#24eb# => X"44004800",
		16#24ec# => X"8681fff8",
		16#24ed# => X"d7e117f0",
		16#24ee# => X"d7e177f4",
		16#24ef# => X"d7e187f8",
		16#24f0# => X"d7e14ffc",
		16#24f1# => X"1a000001",
		16#24f2# => X"9c21ffe0",
		16#24f3# => X"040000a6",
		16#24f4# => X"9dc00000",
		16#24f5# => X"aa10874a",
		16#24f6# => X"a84b0000",
		16#24f7# => X"a880c8ff",
		16#24f8# => X"9dce0001",
		16#24f9# => X"04001022",
		16#24fa# => X"e06e2000",
		16#24fb# => X"18600001",
		16#24fc# => X"d4011000",
		16#24fd# => X"a863872b",
		16#24fe# => X"d4018004",
		16#24ff# => X"d4017008",
		16#2500# => X"0400107e",
		16#2501# => X"d401580c",
		16#2502# => X"bc2e0020",
		16#2503# => X"13fffff5",
		16#2504# => X"a880c8ff",
		16#2505# => X"1a000001",
		16#2506# => X"9dc00000",
		16#2507# => X"aa108754",
		16#2508# => X"a880c93f",
		16#2509# => X"9dce0001",
		16#250a# => X"04001011",
		16#250b# => X"e06e2000",
		16#250c# => X"18600001",
		16#250d# => X"d4011000",
		16#250e# => X"a863872b",
		16#250f# => X"d4018004",
		16#2510# => X"d4017008",
		16#2511# => X"0400106d",
		16#2512# => X"d401580c",
		16#2513# => X"bc2e0020",
		16#2514# => X"13fffff5",
		16#2515# => X"a880c93f",
		16#2516# => X"1a000001",
		16#2517# => X"9dc00000",
		16#2518# => X"aa108617",
		16#2519# => X"a880c9ff",
		16#251a# => X"9dce0001",
		16#251b# => X"04001000",
		16#251c# => X"e06e2000",
		16#251d# => X"18600001",
		16#251e# => X"d4011000",
		16#251f# => X"a863872b",
		16#2520# => X"d4018004",
		16#2521# => X"d4017008",
		16#2522# => X"0400105c",
		16#2523# => X"d401580c",
		16#2524# => X"bc2e0020",
		16#2525# => X"13fffff5",
		16#2526# => X"a880c9ff",
		16#2527# => X"1a000001",
		16#2528# => X"9dc00000",
		16#2529# => X"aa108614",
		16#252a# => X"a880cabf",
		16#252b# => X"9dce0001",
		16#252c# => X"04000fef",
		16#252d# => X"e06e2000",
		16#252e# => X"18600001",
		16#252f# => X"d4011000",
		16#2530# => X"a863872b",
		16#2531# => X"d4018004",
		16#2532# => X"d4017008",
		16#2533# => X"0400104b",
		16#2534# => X"d401580c",
		16#2535# => X"bc2e0020",
		16#2536# => X"13fffff5",
		16#2537# => X"a880cabf",
		16#2538# => X"1a000001",
		16#2539# => X"9dc00000",
		16#253a# => X"aa10861b",
		16#253b# => X"a880caff",
		16#253c# => X"9dce0001",
		16#253d# => X"04000fde",
		16#253e# => X"e06e2000",
		16#253f# => X"18600001",
		16#2540# => X"d4011000",
		16#2541# => X"a863872b",
		16#2542# => X"d4018004",
		16#2543# => X"d4017008",
		16#2544# => X"0400103a",
		16#2545# => X"d401580c",
		16#2546# => X"bc2e0020",
		16#2547# => X"13fffff5",
		16#2548# => X"a880caff",
		16#2549# => X"1a000001",
		16#254a# => X"9dc00000",
		16#254b# => X"aa108622",
		16#254c# => X"a880cb3f",
		16#254d# => X"9dce0001",
		16#254e# => X"04000fcd",
		16#254f# => X"e06e2000",
		16#2550# => X"18600001",
		16#2551# => X"d4011000",
		16#2552# => X"a863872b",
		16#2553# => X"d4018004",
		16#2554# => X"d4017008",
		16#2555# => X"04001029",
		16#2556# => X"d401580c",
		16#2557# => X"bc2e0020",
		16#2558# => X"13fffff5",
		16#2559# => X"a880cb3f",
		16#255a# => X"1a000001",
		16#255b# => X"9dc00000",
		16#255c# => X"aa108629",
		16#255d# => X"a880cb7f",
		16#255e# => X"9dce0001",
		16#255f# => X"04000fbc",
		16#2560# => X"e06e2000",
		16#2561# => X"18600001",
		16#2562# => X"d4011000",
		16#2563# => X"a863872b",
		16#2564# => X"d4018004",
		16#2565# => X"d4017008",
		16#2566# => X"04001018",
		16#2567# => X"d401580c",
		16#2568# => X"bc2e0020",
		16#2569# => X"13fffff5",
		16#256a# => X"a880cb7f",
		16#256b# => X"1a000001",
		16#256c# => X"9dc00000",
		16#256d# => X"aa108630",
		16#256e# => X"a880cbbf",
		16#256f# => X"9dce0001",
		16#2570# => X"04000fab",
		16#2571# => X"e06e2000",
		16#2572# => X"18600001",
		16#2573# => X"d4011000",
		16#2574# => X"a863872b",
		16#2575# => X"d4018004",
		16#2576# => X"d4017008",
		16#2577# => X"04001007",
		16#2578# => X"d401580c",
		16#2579# => X"bc2e0020",
		16#257a# => X"13fffff5",
		16#257b# => X"a880cbbf",
		16#257c# => X"1a000001",
		16#257d# => X"9dc00000",
		16#257e# => X"aa108637",
		16#257f# => X"a880cbff",
		16#2580# => X"9dce0001",
		16#2581# => X"04000f9a",
		16#2582# => X"e06e2000",
		16#2583# => X"18600001",
		16#2584# => X"d4011000",
		16#2585# => X"a863872b",
		16#2586# => X"d4018004",
		16#2587# => X"d4017008",
		16#2588# => X"04000ff6",
		16#2589# => X"d401580c",
		16#258a# => X"bc2e0020",
		16#258b# => X"13fffff5",
		16#258c# => X"a880cbff",
		16#258d# => X"9c210020",
		16#258e# => X"8521fffc",
		16#258f# => X"8441fff0",
		16#2590# => X"85c1fff4",
		16#2591# => X"44004800",
		16#2592# => X"8601fff8",
		16#2593# => X"d7e14ffc",
		16#2594# => X"9c21fffc",
		16#2595# => X"9c210004",
		16#2596# => X"8521fffc",
		16#2597# => X"00000f84",
		16#2598# => X"a860c000",
		16#2599# => X"d7e14ffc",
		16#259a# => X"9c21fffc",
		16#259b# => X"9c210004",
		16#259c# => X"8521fffc",
		16#259d# => X"00000f7e",
		16#259e# => X"a860c002",
		16#259f# => X"9c800001",
		16#25a0# => X"18a00001",
		16#25a1# => X"e0641808",
		16#25a2# => X"a8a5c4b8",
		16#25a3# => X"84850000",
		16#25a4# => X"e0832003",
		16#25a5# => X"bc040000",
		16#25a6# => X"13fffffd",
		16#25a7# => X"15000000",
		16#25a8# => X"44004800",
		16#25a9# => X"15000000",
		16#25aa# => X"18800001",
		16#25ab# => X"9ca00001",
		16#25ac# => X"a884c4b8",
		16#25ad# => X"e0651808",
		16#25ae# => X"84a40000",
		16#25af# => X"e0632804",
		16#25b0# => X"d4041800",
		16#25b1# => X"44004800",
		16#25b2# => X"15000000",
		16#25b3# => X"9ca00001",
		16#25b4# => X"18800001",
		16#25b5# => X"e0651808",
		16#25b6# => X"a884c4b8",
		16#25b7# => X"ac63ffff",
		16#25b8# => X"84a40000",
		16#25b9# => X"e0632803",
		16#25ba# => X"d4041800",
		16#25bb# => X"44004800",
		16#25bc# => X"15000000",
		16#25bd# => X"18600001",
		16#25be# => X"d7e117fc",
		16#25bf# => X"a863c4b8",
		16#25c0# => X"9c400000",
		16#25c1# => X"9c21fffc",
		16#25c2# => X"d4031000",
		16#25c3# => X"9c210004",
		16#25c4# => X"44004800",
		16#25c5# => X"8441fffc",
		16#25c6# => X"18600001",
		16#25c7# => X"9c80ffff",
		16#25c8# => X"a863c4b8",
		16#25c9# => X"d4032000",
		16#25ca# => X"44004800",
		16#25cb# => X"15000000",
		16#25cc# => X"9c21fffc",
		16#25cd# => X"d4014800",
		16#25ce# => X"9d600000",
		16#25cf# => X"9d040000",
		16#25d0# => X"9ca30000",
		16#25d1# => X"e4285800",
		16#25d2# => X"0c000036",
		16#25d3# => X"9ce00000",
		16#25d4# => X"e4482800",
		16#25d5# => X"10000032",
		16#25d6# => X"e4082800",
		16#25d7# => X"1000002e",
		16#25d8# => X"e48b4000",
		16#25d9# => X"0c00000d",
		16#25da# => X"9da00020",
		16#25db# => X"19208000",
		16#25dc# => X"9cc0ffff",
		16#25dd# => X"e0654803",
		16#25de# => X"b8870001",
		16#25df# => X"9de50000",
		16#25e0# => X"b863005f",
		16#25e1# => X"e1ad3000",
		16#25e2# => X"e0e41804",
		16#25e3# => X"e4874000",
		16#25e4# => X"13fffff9",
		16#25e5# => X"b8a50001",
		16#25e6# => X"b8e70041",
		16#25e7# => X"9dad0001",
		16#25e8# => X"9d200000",
		16#25e9# => X"e4896800",
		16#25ea# => X"0c00001e",
		16#25eb# => X"9caf0000",
		16#25ec# => X"19e08000",
		16#25ed# => X"9e200000",
		16#25ee# => X"e0657803",
		16#25ef# => X"b8870001",
		16#25f0# => X"b863005f",
		16#25f1# => X"e0e41804",
		16#25f2# => X"e0c74002",
		16#25f3# => X"e0667803",
		16#25f4# => X"b863005f",
		16#25f5# => X"9c800000",
		16#25f6# => X"e4232000",
		16#25f7# => X"10000003",
		16#25f8# => X"b86b0001",
		16#25f9# => X"9c800001",
		16#25fa# => X"b8a50001",
		16#25fb# => X"e4248800",
		16#25fc# => X"0c000003",
		16#25fd# => X"e1632004",
		16#25fe# => X"9ce60000",
		16#25ff# => X"9d290001",
		16#2600# => X"e4896800",
		16#2601# => X"13ffffed",
		16#2602# => X"15000000",
		16#2603# => X"00000005",
		16#2604# => X"15000000",
		16#2605# => X"00000003",
		16#2606# => X"9d600001",
		16#2607# => X"9ce50000",
		16#2608# => X"85210000",
		16#2609# => X"44004800",
		16#260a# => X"9c210004",
		16#260b# => X"9c21fff8",
		16#260c# => X"d4014800",
		16#260d# => X"d4017004",
		16#260e# => X"9ca30000",
		16#260f# => X"9dc00000",
		16#2610# => X"e5850000",
		16#2611# => X"0c000004",
		16#2612# => X"9c600000",
		16#2613# => X"9dc00001",
		16#2614# => X"e0a02802",
		16#2615# => X"e5840000",
		16#2616# => X"0c000004",
		16#2617# => X"15000000",
		16#2618# => X"9dce0001",
		16#2619# => X"e0802002",
		16#261a# => X"07ffffb2",
		16#261b# => X"9c650000",
		16#261c# => X"bc0e0001",
		16#261d# => X"0c000003",
		16#261e# => X"15000000",
		16#261f# => X"e1605802",
		16#2620# => X"85210000",
		16#2621# => X"85c10004",
		16#2622# => X"44004800",
		16#2623# => X"9c210008",
		16#2624# => X"d7e117f8",
		16#2625# => X"18400001",
		16#2626# => X"d7e14ffc",
		16#2627# => X"a8428760",
		16#2628# => X"9c21fff0",
		16#2629# => X"84a20000",
		16#262a# => X"84c20004",
		16#262b# => X"d4011800",
		16#262c# => X"d4012004",
		16#262d# => X"0400094c",
		16#262e# => X"15000000",
		16#262f# => X"bd6b0000",
		16#2630# => X"1000000a",
		16#2631# => X"15000000",
		16#2632# => X"84610000",
		16#2633# => X"84810004",
		16#2634# => X"04000a40",
		16#2635# => X"15000000",
		16#2636# => X"9c210010",
		16#2637# => X"8521fffc",
		16#2638# => X"44004800",
		16#2639# => X"8441fff8",
		16#263a# => X"84a20000",
		16#263b# => X"84c20004",
		16#263c# => X"84610000",
		16#263d# => X"84810004",
		16#263e# => X"040006a9",
		16#263f# => X"18408000",
		16#2640# => X"e06b0004",
		16#2641# => X"e08c0004",
		16#2642# => X"04000a32",
		16#2643# => X"15000000",
		16#2644# => X"9c210010",
		16#2645# => X"8521fffc",
		16#2646# => X"e16b1000",
		16#2647# => X"44004800",
		16#2648# => X"8441fff8",
		16#2649# => X"d7e117fc",
		16#264a# => X"84c30000",
		16#264b# => X"bca60001",
		16#264c# => X"1000004e",
		16#264d# => X"9c21fffc",
		16#264e# => X"84e40000",
		16#264f# => X"bca70001",
		16#2650# => X"1000006e",
		16#2651# => X"bc260004",
		16#2652# => X"0c000083",
		16#2653# => X"bc070004",
		16#2654# => X"1000006a",
		16#2655# => X"bc270002",
		16#2656# => X"0c000055",
		16#2657# => X"bc060002",
		16#2658# => X"10000066",
		16#2659# => X"15000000",
		16#265a# => X"84e30008",
		16#265b# => X"85a40008",
		16#265c# => X"8583000c",
		16#265d# => X"e1676802",
		16#265e# => X"b9eb009f",
		16#265f# => X"e0cf5805",
		16#2660# => X"e0c67802",
		16#2661# => X"bd46001f",
		16#2662# => X"1000003c",
		16#2663# => X"8504000c",
		16#2664# => X"bdab0000",
		16#2665# => X"10000064",
		16#2666# => X"9da00001",
		16#2667# => X"e1683048",
		16#2668# => X"e0cd3008",
		16#2669# => X"9cc6ffff",
		16#266a# => X"e1064003",
		16#266b# => X"e0c04002",
		16#266c# => X"e1064004",
		16#266d# => X"b908005f",
		16#266e# => X"e1085804",
		16#266f# => X"84630004",
		16#2670# => X"84840004",
		16#2671# => X"e4032000",
		16#2672# => X"10000035",
		16#2673# => X"e0886000",
		16#2674# => X"bc030000",
		16#2675# => X"10000003",
		16#2676# => X"e08c4002",
		16#2677# => X"e0886002",
		16#2678# => X"bd840000",
		16#2679# => X"1000004a",
		16#267a# => X"9c400000",
		16#267b# => X"d4053808",
		16#267c# => X"d4051004",
		16#267d# => X"d405200c",
		16#267e# => X"18403fff",
		16#267f# => X"9c64ffff",
		16#2680# => X"a842fffe",
		16#2681# => X"e4431000",
		16#2682# => X"1000000d",
		16#2683# => X"9cc00003",
		16#2684# => X"84650008",
		16#2685# => X"e0842000",
		16#2686# => X"18403fff",
		16#2687# => X"9cc4ffff",
		16#2688# => X"a842fffe",
		16#2689# => X"e4a61000",
		16#268a# => X"13fffffb",
		16#268b# => X"9c63ffff",
		16#268c# => X"d405200c",
		16#268d# => X"d4051808",
		16#268e# => X"9cc00003",
		16#268f# => X"a8650000",
		16#2690# => X"bd640000",
		16#2691# => X"10000009",
		16#2692# => X"d4053000",
		16#2693# => X"b8c40041",
		16#2694# => X"84a50008",
		16#2695# => X"a4840001",
		16#2696# => X"9ca50001",
		16#2697# => X"e0843004",
		16#2698# => X"d4032808",
		16#2699# => X"d403200c",
		16#269a# => X"9c210004",
		16#269b# => X"a9630000",
		16#269c# => X"44004800",
		16#269d# => X"8441fffc",
		16#269e# => X"e5a76800",
		16#269f# => X"1000001c",
		16#26a0# => X"15000000",
		16#26a1# => X"84630004",
		16#26a2# => X"84840004",
		16#26a3# => X"e4032000",
		16#26a4# => X"0fffffd0",
		16#26a5# => X"9d000000",
		16#26a6# => X"e0886000",
		16#26a7# => X"d4051804",
		16#26a8# => X"d4053808",
		16#26a9# => X"03ffffe5",
		16#26aa# => X"d405200c",
		16#26ab# => X"bc260002",
		16#26ac# => X"13ffffee",
		16#26ad# => X"15000000",
		16#26ae# => X"d4053000",
		16#26af# => X"84c30004",
		16#26b0# => X"d4053004",
		16#26b1# => X"84c30008",
		16#26b2# => X"d4053008",
		16#26b3# => X"84c3000c",
		16#26b4# => X"d405300c",
		16#26b5# => X"84c30004",
		16#26b6# => X"84840004",
		16#26b7# => X"a8650000",
		16#26b8# => X"e0843003",
		16#26b9# => X"03ffffe1",
		16#26ba# => X"d4052004",
		16#26bb# => X"a8ed0000",
		16#26bc# => X"03ffffb3",
		16#26bd# => X"9d800000",
		16#26be# => X"a8640000",
		16#26bf# => X"9c210004",
		16#26c0# => X"a9630000",
		16#26c1# => X"44004800",
		16#26c2# => X"8441fffc",
		16#26c3# => X"e0802002",
		16#26c4# => X"9c600001",
		16#26c5# => X"d4053808",
		16#26c6# => X"d4051804",
		16#26c7# => X"03ffffb7",
		16#26c8# => X"d405200c",
		16#26c9# => X"bc0b0000",
		16#26ca# => X"13ffffa5",
		16#26cb# => X"e16c3048",
		16#26cc# => X"e1ad3008",
		16#26cd# => X"e0e73000",
		16#26ce# => X"9ccdffff",
		16#26cf# => X"e1866003",
		16#26d0# => X"e0c06002",
		16#26d1# => X"e1866004",
		16#26d2# => X"b98c005f",
		16#26d3# => X"03ffff9c",
		16#26d4# => X"e18c5804",
		16#26d5# => X"bc270004",
		16#26d6# => X"13ffffc4",
		16#26d7# => X"15000000",
		16#26d8# => X"84a30004",
		16#26d9# => X"84840004",
		16#26da# => X"e4252000",
		16#26db# => X"0fffffbf",
		16#26dc# => X"15000000",
		16#26dd# => X"18600001",
		16#26de# => X"03ffffbc",
		16#26df# => X"a863876c",
		16#26e0# => X"d7e117fc",
		16#26e1# => X"84a30000",
		16#26e2# => X"9c21fffc",
		16#26e3# => X"8483000c",
		16#26e4# => X"bc450001",
		16#26e5# => X"0c00003d",
		16#26e6# => X"84c30004",
		16#26e7# => X"bc050004",
		16#26e8# => X"10000037",
		16#26e9# => X"bc050002",
		16#26ea# => X"10000024",
		16#26eb# => X"bc040000",
		16#26ec# => X"1000001b",
		16#26ed# => X"15000000",
		16#26ee# => X"84630008",
		16#26ef# => X"bd63ff82",
		16#26f0# => X"0c000039",
		16#26f1# => X"bd43007f",
		16#26f2# => X"1000002d",
		16#26f3# => X"a4a4007f",
		16#26f4# => X"bc250040",
		16#26f5# => X"0c000021",
		16#26f6# => X"9c63007f",
		16#26f7# => X"9c84003f",
		16#26f8# => X"bd640000",
		16#26f9# => X"0c000023",
		16#26fa# => X"15000000",
		16#26fb# => X"1840007f",
		16#26fc# => X"b8a40047",
		16#26fd# => X"a842ffff",
		16#26fe# => X"a48300ff",
		16#26ff# => X"e0651003",
		16#2700# => X"b8840017",
		16#2701# => X"b8a6001f",
		16#2702# => X"e0832004",
		16#2703# => X"9c210004",
		16#2704# => X"e1642804",
		16#2705# => X"44004800",
		16#2706# => X"8441fffc",
		16#2707# => X"a8640000",
		16#2708# => X"b8a6001f",
		16#2709# => X"e0832004",
		16#270a# => X"9c210004",
		16#270b# => X"e1642804",
		16#270c# => X"44004800",
		16#270d# => X"8441fffc",
		16#270e# => X"9c800000",
		16#270f# => X"b8a6001f",
		16#2710# => X"a8640000",
		16#2711# => X"9c210004",
		16#2712# => X"e0832004",
		16#2713# => X"8441fffc",
		16#2714# => X"44004800",
		16#2715# => X"e1642804",
		16#2716# => X"a4a40080",
		16#2717# => X"bc050000",
		16#2718# => X"13ffffe1",
		16#2719# => X"bd640000",
		16#271a# => X"03ffffde",
		16#271b# => X"9c840040",
		16#271c# => X"b8840041",
		16#271d# => X"03ffffde",
		16#271e# => X"9c630001",
		16#271f# => X"18807f80",
		16#2720# => X"03ffffe1",
		16#2721# => X"9c600000",
		16#2722# => X"18400010",
		16#2723# => X"e0641004",
		16#2724# => X"1840007f",
		16#2725# => X"18807f80",
		16#2726# => X"a842ffff",
		16#2727# => X"03ffffda",
		16#2728# => X"e0631003",
		16#2729# => X"9ce0ff82",
		16#272a# => X"e0671802",
		16#272b# => X"bd430019",
		16#272c# => X"1000001f",
		16#272d# => X"9ca00000",
		16#272e# => X"9ce00001",
		16#272f# => X"e0a41848",
		16#2730# => X"e0671808",
		16#2731# => X"9c63ffff",
		16#2732# => X"e0832003",
		16#2733# => X"e0602002",
		16#2734# => X"e0632004",
		16#2735# => X"b863005f",
		16#2736# => X"e0a32804",
		16#2737# => X"a465007f",
		16#2738# => X"bc230040",
		16#2739# => X"10000012",
		16#273a# => X"15000000",
		16#273b# => X"a4650080",
		16#273c# => X"bc030000",
		16#273d# => X"10000004",
		16#273e# => X"18403fff",
		16#273f# => X"9ca50040",
		16#2740# => X"18403fff",
		16#2741# => X"b8650047",
		16#2742# => X"a842ffff",
		16#2743# => X"9c800001",
		16#2744# => X"e4451000",
		16#2745# => X"1840007f",
		16#2746# => X"a842ffff",
		16#2747# => X"13ffffb9",
		16#2748# => X"e0631003",
		16#2749# => X"03ffffb7",
		16#274a# => X"9c800000",
		16#274b# => X"03fffff5",
		16#274c# => X"9ca5003f",
		16#274d# => X"d7e117fc",
		16#274e# => X"1840007f",
		16#274f# => X"84a30000",
		16#2750# => X"a842ffff",
		16#2751# => X"b8c50057",
		16#2752# => X"b8e5005f",
		16#2753# => X"9c21fffc",
		16#2754# => X"a4c600ff",
		16#2755# => X"d4043804",
		16#2756# => X"bc260000",
		16#2757# => X"10000016",
		16#2758# => X"e0651003",
		16#2759# => X"bc230000",
		16#275a# => X"0c000020",
		16#275b# => X"9ca0ff82",
		16#275c# => X"b8630007",
		16#275d# => X"d4042808",
		16#275e# => X"9ca00003",
		16#275f# => X"d4042800",
		16#2760# => X"9ca0ff81",
		16#2761# => X"18403fff",
		16#2762# => X"e0631800",
		16#2763# => X"a842ffff",
		16#2764# => X"a8c50000",
		16#2765# => X"e4a31000",
		16#2766# => X"13fffffb",
		16#2767# => X"9ca5ffff",
		16#2768# => X"9c210004",
		16#2769# => X"d4043008",
		16#276a# => X"d404180c",
		16#276b# => X"44004800",
		16#276c# => X"8441fffc",
		16#276d# => X"bc2600ff",
		16#276e# => X"0c000011",
		16#276f# => X"9cc6ff81",
		16#2770# => X"b8630007",
		16#2771# => X"18404000",
		16#2772# => X"d4043008",
		16#2773# => X"e0631004",
		16#2774# => X"9ca00003",
		16#2775# => X"d4042800",
		16#2776# => X"d404180c",
		16#2777# => X"9c210004",
		16#2778# => X"44004800",
		16#2779# => X"8441fffc",
		16#277a# => X"9c600002",
		16#277b# => X"9c210004",
		16#277c# => X"d4041800",
		16#277d# => X"44004800",
		16#277e# => X"8441fffc",
		16#277f# => X"bc230000",
		16#2780# => X"0c00000a",
		16#2781# => X"15000000",
		16#2782# => X"18400010",
		16#2783# => X"e0a51003",
		16#2784# => X"bc050000",
		16#2785# => X"13fffff0",
		16#2786# => X"15000000",
		16#2787# => X"9ca00001",
		16#2788# => X"03ffffee",
		16#2789# => X"d4042800",
		16#278a# => X"9c600004",
		16#278b# => X"03ffffec",
		16#278c# => X"d4041800",
		16#278d# => X"d7e14ffc",
		16#278e# => X"d7e117f4",
		16#278f# => X"d7e177f8",
		16#2790# => X"9c21ffbc",
		16#2791# => X"9dc10020",
		16#2792# => X"d4011834",
		16#2793# => X"d4012030",
		16#2794# => X"9c610034",
		16#2795# => X"a88e0000",
		16#2796# => X"07ffffb7",
		16#2797# => X"9c410010",
		16#2798# => X"9c610030",
		16#2799# => X"07ffffb4",
		16#279a# => X"a8820000",
		16#279b# => X"a86e0000",
		16#279c# => X"a8820000",
		16#279d# => X"07fffeac",
		16#279e# => X"a8a10000",
		16#279f# => X"07ffff41",
		16#27a0# => X"a86b0000",
		16#27a1# => X"9c210044",
		16#27a2# => X"8521fffc",
		16#27a3# => X"8441fff4",
		16#27a4# => X"44004800",
		16#27a5# => X"85c1fff8",
		16#27a6# => X"d7e14ffc",
		16#27a7# => X"d7e117f4",
		16#27a8# => X"d7e177f8",
		16#27a9# => X"9c21ffbc",
		16#27aa# => X"9dc10020",
		16#27ab# => X"d4011834",
		16#27ac# => X"d4012030",
		16#27ad# => X"9c610034",
		16#27ae# => X"a88e0000",
		16#27af# => X"07ffff9e",
		16#27b0# => X"9c410010",
		16#27b1# => X"9c610030",
		16#27b2# => X"07ffff9b",
		16#27b3# => X"a8820000",
		16#27b4# => X"84c10014",
		16#27b5# => X"a86e0000",
		16#27b6# => X"acc60001",
		16#27b7# => X"a8820000",
		16#27b8# => X"a8a10000",
		16#27b9# => X"07fffe90",
		16#27ba# => X"d4013014",
		16#27bb# => X"07ffff25",
		16#27bc# => X"a86b0000",
		16#27bd# => X"9c210044",
		16#27be# => X"8521fffc",
		16#27bf# => X"8441fff4",
		16#27c0# => X"44004800",
		16#27c1# => X"85c1fff8",
		16#27c2# => X"d7e14ffc",
		16#27c3# => X"d7e117f4",
		16#27c4# => X"d7e177f8",
		16#27c5# => X"9c21ffbc",
		16#27c6# => X"9c410020",
		16#27c7# => X"d4011834",
		16#27c8# => X"d4012030",
		16#27c9# => X"9c610034",
		16#27ca# => X"a8820000",
		16#27cb# => X"07ffff82",
		16#27cc# => X"9dc10010",
		16#27cd# => X"9c610030",
		16#27ce# => X"07ffff7f",
		16#27cf# => X"a88e0000",
		16#27d0# => X"84a10020",
		16#27d1# => X"bc450001",
		16#27d2# => X"0c00005e",
		16#27d3# => X"84c10010",
		16#27d4# => X"bc460001",
		16#27d5# => X"0c00006d",
		16#27d6# => X"bc250004",
		16#27d7# => X"0c000055",
		16#27d8# => X"bc260004",
		16#27d9# => X"0c000065",
		16#27da# => X"bc250002",
		16#27db# => X"0c000055",
		16#27dc# => X"bc260002",
		16#27dd# => X"0c000065",
		16#27de# => X"9c600000",
		16#27df# => X"8481001c",
		16#27e0# => X"a8a30000",
		16#27e1# => X"04000916",
		16#27e2# => X"84c1002c",
		16#27e3# => X"84610024",
		16#27e4# => X"84410014",
		16#27e5# => X"84810028",
		16#27e6# => X"e0431005",
		16#27e7# => X"84a10018",
		16#27e8# => X"e0601002",
		16#27e9# => X"e0852000",
		16#27ea# => X"e0431004",
		16#27eb# => X"9c640002",
		16#27ec# => X"b842005f",
		16#27ed# => X"d4011808",
		16#27ee# => X"bd6b0000",
		16#27ef# => X"d4011004",
		16#27f0# => X"10000008",
		16#27f1# => X"a86b0000",
		16#27f2# => X"a44b0001",
		16#27f3# => X"bc020000",
		16#27f4# => X"0c00002a",
		16#27f5# => X"9c840003",
		16#27f6# => X"b86b0041",
		16#27f7# => X"d4012008",
		16#27f8# => X"18403fff",
		16#27f9# => X"a842ffff",
		16#27fa# => X"e4431000",
		16#27fb# => X"10000014",
		16#27fc# => X"84810008",
		16#27fd# => X"00000008",
		16#27fe# => X"e0631800",
		16#27ff# => X"18403fff",
		16#2800# => X"a842ffff",
		16#2801# => X"e4a31000",
		16#2802# => X"0c00000c",
		16#2803# => X"e18c6000",
		16#2804# => X"e0631800",
		16#2805# => X"bd6c0000",
		16#2806# => X"13fffff9",
		16#2807# => X"9c84ffff",
		16#2808# => X"18403fff",
		16#2809# => X"a8630001",
		16#280a# => X"a842ffff",
		16#280b# => X"e4a31000",
		16#280c# => X"13fffff8",
		16#280d# => X"e18c6000",
		16#280e# => X"d4012008",
		16#280f# => X"a443007f",
		16#2810# => X"bc220040",
		16#2811# => X"0c000011",
		16#2812# => X"a4430080",
		16#2813# => X"9c400003",
		16#2814# => X"d401180c",
		16#2815# => X"d4011000",
		16#2816# => X"a8610000",
		16#2817# => X"07fffec9",
		16#2818# => X"15000000",
		16#2819# => X"9c210044",
		16#281a# => X"8521fffc",
		16#281b# => X"8441fff4",
		16#281c# => X"44004800",
		16#281d# => X"85c1fff8",
		16#281e# => X"b98c0041",
		16#281f# => X"18408000",
		16#2820# => X"03ffffd6",
		16#2821# => X"e18c1004",
		16#2822# => X"bc220000",
		16#2823# => X"13fffff1",
		16#2824# => X"9c400003",
		16#2825# => X"bc0c0000",
		16#2826# => X"13ffffee",
		16#2827# => X"15000000",
		16#2828# => X"9c630040",
		16#2829# => X"9c40ff80",
		16#282a# => X"03ffffe9",
		16#282b# => X"e0631003",
		16#282c# => X"18600001",
		16#282d# => X"bc060002",
		16#282e# => X"13ffffe9",
		16#282f# => X"a863876c",
		16#2830# => X"84810024",
		16#2831# => X"a8620000",
		16#2832# => X"84410014",
		16#2833# => X"e0441005",
		16#2834# => X"e0801002",
		16#2835# => X"e0441004",
		16#2836# => X"b842005f",
		16#2837# => X"07fffea9",
		16#2838# => X"d4011024",
		16#2839# => X"9c210044",
		16#283a# => X"8521fffc",
		16#283b# => X"8441fff4",
		16#283c# => X"44004800",
		16#283d# => X"85c1fff8",
		16#283e# => X"18600001",
		16#283f# => X"bc050002",
		16#2840# => X"13ffffd7",
		16#2841# => X"a863876c",
		16#2842# => X"84410014",
		16#2843# => X"84810024",
		16#2844# => X"a86e0000",
		16#2845# => X"e0441005",
		16#2846# => X"e0801002",
		16#2847# => X"e0441004",
		16#2848# => X"b842005f",
		16#2849# => X"07fffe97",
		16#284a# => X"d4011014",
		16#284b# => X"9c210044",
		16#284c# => X"8521fffc",
		16#284d# => X"8441fff4",
		16#284e# => X"44004800",
		16#284f# => X"85c1fff8",
		16#2850# => X"d7e14ffc",
		16#2851# => X"d7e117f4",
		16#2852# => X"d7e177f8",
		16#2853# => X"9c21ffcc",
		16#2854# => X"9c410010",
		16#2855# => X"d4011824",
		16#2856# => X"d4012020",
		16#2857# => X"9c610024",
		16#2858# => X"07fffef5",
		16#2859# => X"a8820000",
		16#285a# => X"9c610020",
		16#285b# => X"07fffef2",
		16#285c# => X"a8810000",
		16#285d# => X"84a10010",
		16#285e# => X"bca50001",
		16#285f# => X"1000002c",
		16#2860# => X"a8620000",
		16#2861# => X"84c10000",
		16#2862# => X"bca60001",
		16#2863# => X"10000028",
		16#2864# => X"a8610000",
		16#2865# => X"84810014",
		16#2866# => X"84610004",
		16#2867# => X"bc050004",
		16#2868# => X"e0641805",
		16#2869# => X"1000002d",
		16#286a# => X"d4011814",
		16#286b# => X"bc250002",
		16#286c# => X"0c00002a",
		16#286d# => X"bc260004",
		16#286e# => X"0c000040",
		16#286f# => X"bc260002",
		16#2870# => X"0c000035",
		16#2871# => X"84a10018",
		16#2872# => X"84810008",
		16#2873# => X"8461001c",
		16#2874# => X"e0852002",
		16#2875# => X"84e1000c",
		16#2876# => X"e4633800",
		16#2877# => X"0c00001b",
		16#2878# => X"d4012018",
		16#2879# => X"9ca0001f",
		16#287a# => X"18c04000",
		16#287b# => X"9d000000",
		16#287c# => X"e4471800",
		16#287d# => X"10000004",
		16#287e# => X"9ca5ffff",
		16#287f# => X"e1083004",
		16#2880# => X"e0633802",
		16#2881# => X"b8c60041",
		16#2882# => X"bc250000",
		16#2883# => X"13fffff9",
		16#2884# => X"e0631800",
		16#2885# => X"a488007f",
		16#2886# => X"bc240040",
		16#2887# => X"0c000015",
		16#2888# => X"a4880080",
		16#2889# => X"d401401c",
		16#288a# => X"a8620000",
		16#288b# => X"07fffe55",
		16#288c# => X"15000000",
		16#288d# => X"9c210034",
		16#288e# => X"8521fffc",
		16#288f# => X"8441fff4",
		16#2890# => X"44004800",
		16#2891# => X"85c1fff8",
		16#2892# => X"9c84ffff",
		16#2893# => X"e0631800",
		16#2894# => X"03ffffe5",
		16#2895# => X"d4012018",
		16#2896# => X"18600001",
		16#2897# => X"e4053000",
		16#2898# => X"0ffffff2",
		16#2899# => X"a863876c",
		16#289a# => X"03fffff1",
		16#289b# => X"15000000",
		16#289c# => X"bc240000",
		16#289d# => X"13ffffec",
		16#289e# => X"bc030000",
		16#289f# => X"13ffffea",
		16#28a0# => X"9c60ff80",
		16#28a1# => X"9d080040",
		16#28a2# => X"e1081803",
		16#28a3# => X"03ffffe7",
		16#28a4# => X"d401401c",
		16#28a5# => X"a8620000",
		16#28a6# => X"9c400004",
		16#28a7# => X"07fffe39",
		16#28a8# => X"d4011010",
		16#28a9# => X"9c210034",
		16#28aa# => X"8521fffc",
		16#28ab# => X"8441fff4",
		16#28ac# => X"44004800",
		16#28ad# => X"85c1fff8",
		16#28ae# => X"9c600000",
		16#28af# => X"d401181c",
		16#28b0# => X"d4011818",
		16#28b1# => X"03ffffda",
		16#28b2# => X"a8620000",
		16#28b3# => X"84a30000",
		16#28b4# => X"9d600001",
		16#28b5# => X"e4a55800",
		16#28b6# => X"10000016",
		16#28b7# => X"15000000",
		16#28b8# => X"84c40000",
		16#28b9# => X"e4a65800",
		16#28ba# => X"10000012",
		16#28bb# => X"bc250004",
		16#28bc# => X"0c000037",
		16#28bd# => X"bc260004",
		16#28be# => X"0c000019",
		16#28bf# => X"bc250002",
		16#28c0# => X"0c000014",
		16#28c1# => X"bc260002",
		16#28c2# => X"0c00000c",
		16#28c3# => X"15000000",
		16#28c4# => X"84a30004",
		16#28c5# => X"84c40004",
		16#28c6# => X"e4053000",
		16#28c7# => X"10000016",
		16#28c8# => X"15000000",
		16#28c9# => X"bc050000",
		16#28ca# => X"0c000008",
		16#28cb# => X"15000000",
		16#28cc# => X"44004800",
		16#28cd# => X"15000000",
		16#28ce# => X"84630004",
		16#28cf# => X"bc030000",
		16#28d0# => X"13fffffc",
		16#28d1# => X"15000000",
		16#28d2# => X"44004800",
		16#28d3# => X"9d60ffff",
		16#28d4# => X"bc060002",
		16#28d5# => X"13fffff7",
		16#28d6# => X"9d600000",
		16#28d7# => X"84640004",
		16#28d8# => X"bc030000",
		16#28d9# => X"13fffff3",
		16#28da# => X"9d60ffff",
		16#28db# => X"44004800",
		16#28dc# => X"9d600001",
		16#28dd# => X"84e30008",
		16#28de# => X"84c40008",
		16#28df# => X"e5a73000",
		16#28e0# => X"0fffffea",
		16#28e1# => X"bc050000",
		16#28e2# => X"e5673000",
		16#28e3# => X"0c00000c",
		16#28e4# => X"bc050000",
		16#28e5# => X"84c3000c",
		16#28e6# => X"8464000c",
		16#28e7# => X"e4a61800",
		16#28e8# => X"10000004",
		16#28e9# => X"e4661800",
		16#28ea# => X"03ffffdf",
		16#28eb# => X"9d600001",
		16#28ec# => X"13ffffe0",
		16#28ed# => X"9d600000",
		16#28ee# => X"bc050000",
		16#28ef# => X"0fffffec",
		16#28f0# => X"9d60ffff",
		16#28f1# => X"44004800",
		16#28f2# => X"15000000",
		16#28f3# => X"13ffffdb",
		16#28f4# => X"15000000",
		16#28f5# => X"85640004",
		16#28f6# => X"84630004",
		16#28f7# => X"44004800",
		16#28f8# => X"e16b1802",
		16#28f9# => X"d7e14ffc",
		16#28fa# => X"d7e117f4",
		16#28fb# => X"d7e177f8",
		16#28fc# => X"9c21ffcc",
		16#28fd# => X"9dc10010",
		16#28fe# => X"d4011824",
		16#28ff# => X"d4012020",
		16#2900# => X"9c610024",
		16#2901# => X"07fffe4c",
		16#2902# => X"a88e0000",
		16#2903# => X"9c610020",
		16#2904# => X"07fffe49",
		16#2905# => X"a8810000",
		16#2906# => X"a86e0000",
		16#2907# => X"07ffffac",
		16#2908# => X"a8810000",
		16#2909# => X"9c210034",
		16#290a# => X"8521fffc",
		16#290b# => X"8441fff4",
		16#290c# => X"44004800",
		16#290d# => X"85c1fff8",
		16#290e# => X"d7e14ffc",
		16#290f# => X"d7e177f8",
		16#2910# => X"d7e117f4",
		16#2911# => X"9c21ffcc",
		16#2912# => X"9dc10010",
		16#2913# => X"d4011824",
		16#2914# => X"d4012020",
		16#2915# => X"9c610024",
		16#2916# => X"07fffe37",
		16#2917# => X"a88e0000",
		16#2918# => X"9c610020",
		16#2919# => X"07fffe34",
		16#291a# => X"a8810000",
		16#291b# => X"9d600001",
		16#291c# => X"84610010",
		16#291d# => X"e4a35800",
		16#291e# => X"10000007",
		16#291f# => X"84610000",
		16#2920# => X"e4a35800",
		16#2921# => X"10000004",
		16#2922# => X"a86e0000",
		16#2923# => X"07ffff90",
		16#2924# => X"a8810000",
		16#2925# => X"9c210034",
		16#2926# => X"8521fffc",
		16#2927# => X"8441fff4",
		16#2928# => X"44004800",
		16#2929# => X"85c1fff8",
		16#292a# => X"d7e14ffc",
		16#292b# => X"d7e177f8",
		16#292c# => X"d7e117f4",
		16#292d# => X"9c21ffcc",
		16#292e# => X"9dc10010",
		16#292f# => X"d4011824",
		16#2930# => X"d4012020",
		16#2931# => X"9c610024",
		16#2932# => X"07fffe1b",
		16#2933# => X"a88e0000",
		16#2934# => X"9c610020",
		16#2935# => X"07fffe18",
		16#2936# => X"a8810000",
		16#2937# => X"9d600001",
		16#2938# => X"84610010",
		16#2939# => X"e4a35800",
		16#293a# => X"10000007",
		16#293b# => X"84610000",
		16#293c# => X"e4a35800",
		16#293d# => X"10000004",
		16#293e# => X"a86e0000",
		16#293f# => X"07ffff74",
		16#2940# => X"a8810000",
		16#2941# => X"9c210034",
		16#2942# => X"8521fffc",
		16#2943# => X"8441fff4",
		16#2944# => X"44004800",
		16#2945# => X"85c1fff8",
		16#2946# => X"d7e14ffc",
		16#2947# => X"d7e177f8",
		16#2948# => X"d7e117f4",
		16#2949# => X"9c21ffcc",
		16#294a# => X"9dc10010",
		16#294b# => X"d4011824",
		16#294c# => X"d4012020",
		16#294d# => X"9c610024",
		16#294e# => X"07fffdff",
		16#294f# => X"a88e0000",
		16#2950# => X"9c610020",
		16#2951# => X"07fffdfc",
		16#2952# => X"a8810000",
		16#2953# => X"84610010",
		16#2954# => X"bca30001",
		16#2955# => X"10000008",
		16#2956# => X"9d60ffff",
		16#2957# => X"84610000",
		16#2958# => X"bca30001",
		16#2959# => X"10000004",
		16#295a# => X"a86e0000",
		16#295b# => X"07ffff58",
		16#295c# => X"a8810000",
		16#295d# => X"9c210034",
		16#295e# => X"8521fffc",
		16#295f# => X"8441fff4",
		16#2960# => X"44004800",
		16#2961# => X"85c1fff8",
		16#2962# => X"d7e14ffc",
		16#2963# => X"d7e177f8",
		16#2964# => X"d7e117f4",
		16#2965# => X"9c21ffcc",
		16#2966# => X"9dc10010",
		16#2967# => X"d4011824",
		16#2968# => X"d4012020",
		16#2969# => X"9c610024",
		16#296a# => X"07fffde3",
		16#296b# => X"a88e0000",
		16#296c# => X"9c610020",
		16#296d# => X"07fffde0",
		16#296e# => X"a8810000",
		16#296f# => X"84610010",
		16#2970# => X"bca30001",
		16#2971# => X"10000008",
		16#2972# => X"9d60ffff",
		16#2973# => X"84610000",
		16#2974# => X"bca30001",
		16#2975# => X"10000004",
		16#2976# => X"a86e0000",
		16#2977# => X"07ffff3c",
		16#2978# => X"a8810000",
		16#2979# => X"9c210034",
		16#297a# => X"8521fffc",
		16#297b# => X"8441fff4",
		16#297c# => X"44004800",
		16#297d# => X"85c1fff8",
		16#297e# => X"d7e14ffc",
		16#297f# => X"d7e177f8",
		16#2980# => X"d7e117f4",
		16#2981# => X"9c21ffcc",
		16#2982# => X"9dc10010",
		16#2983# => X"d4011824",
		16#2984# => X"d4012020",
		16#2985# => X"9c610024",
		16#2986# => X"07fffdc7",
		16#2987# => X"a88e0000",
		16#2988# => X"9c610020",
		16#2989# => X"07fffdc4",
		16#298a# => X"a8810000",
		16#298b# => X"9d600001",
		16#298c# => X"84610010",
		16#298d# => X"e4a35800",
		16#298e# => X"10000007",
		16#298f# => X"84610000",
		16#2990# => X"e4a35800",
		16#2991# => X"10000004",
		16#2992# => X"a86e0000",
		16#2993# => X"07ffff20",
		16#2994# => X"a8810000",
		16#2995# => X"9c210034",
		16#2996# => X"8521fffc",
		16#2997# => X"8441fff4",
		16#2998# => X"44004800",
		16#2999# => X"85c1fff8",
		16#299a# => X"d7e14ffc",
		16#299b# => X"d7e177f8",
		16#299c# => X"d7e117f4",
		16#299d# => X"9c21ffcc",
		16#299e# => X"9dc10010",
		16#299f# => X"d4011824",
		16#29a0# => X"d4012020",
		16#29a1# => X"9c610024",
		16#29a2# => X"07fffdab",
		16#29a3# => X"a88e0000",
		16#29a4# => X"9c610020",
		16#29a5# => X"07fffda8",
		16#29a6# => X"a8810000",
		16#29a7# => X"9d600001",
		16#29a8# => X"84610010",
		16#29a9# => X"e4a35800",
		16#29aa# => X"10000007",
		16#29ab# => X"84610000",
		16#29ac# => X"e4a35800",
		16#29ad# => X"10000004",
		16#29ae# => X"a86e0000",
		16#29af# => X"07ffff04",
		16#29b0# => X"a8810000",
		16#29b1# => X"9c210034",
		16#29b2# => X"8521fffc",
		16#29b3# => X"8441fff4",
		16#29b4# => X"44004800",
		16#29b5# => X"85c1fff8",
		16#29b6# => X"d7e14ffc",
		16#29b7# => X"9c21ffd4",
		16#29b8# => X"d4011824",
		16#29b9# => X"d4012020",
		16#29ba# => X"9c610024",
		16#29bb# => X"07fffd92",
		16#29bc# => X"9c810010",
		16#29bd# => X"9c610020",
		16#29be# => X"07fffd8f",
		16#29bf# => X"a8810000",
		16#29c0# => X"9d600001",
		16#29c1# => X"84610010",
		16#29c2# => X"e4a35800",
		16#29c3# => X"10000005",
		16#29c4# => X"84610000",
		16#29c5# => X"e4a35800",
		16#29c6# => X"0c000006",
		16#29c7# => X"15000000",
		16#29c8# => X"9c21002c",
		16#29c9# => X"8521fffc",
		16#29ca# => X"44004800",
		16#29cb# => X"15000000",
		16#29cc# => X"9c21002c",
		16#29cd# => X"8521fffc",
		16#29ce# => X"44004800",
		16#29cf# => X"9d600000",
		16#29d0# => X"b883005f",
		16#29d1# => X"d7e117f8",
		16#29d2# => X"d7e14ffc",
		16#29d3# => X"9c400003",
		16#29d4# => X"9c21ffe8",
		16#29d5# => X"bc230000",
		16#29d6# => X"d4011000",
		16#29d7# => X"1000000a",
		16#29d8# => X"d4012004",
		16#29d9# => X"9c400002",
		16#29da# => X"d4011000",
		16#29db# => X"07fffd05",
		16#29dc# => X"a8610000",
		16#29dd# => X"9c210018",
		16#29de# => X"8521fffc",
		16#29df# => X"44004800",
		16#29e0# => X"8441fff8",
		16#29e1# => X"a8430000",
		16#29e2# => X"9c60001e",
		16#29e3# => X"bc040000",
		16#29e4# => X"10000007",
		16#29e5# => X"d4011808",
		16#29e6# => X"18608000",
		16#29e7# => X"e4021800",
		16#29e8# => X"1000000f",
		16#29e9# => X"15000000",
		16#29ea# => X"e0401002",
		16#29eb# => X"a8620000",
		16#29ec# => X"04000750",
		16#29ed# => X"d401100c",
		16#29ee# => X"9d6bffff",
		16#29ef# => X"bdab0000",
		16#29f0# => X"13ffffeb",
		16#29f1# => X"9c60001e",
		16#29f2# => X"e0425808",
		16#29f3# => X"e1635802",
		16#29f4# => X"d401100c",
		16#29f5# => X"03ffffe6",
		16#29f6# => X"d4015808",
		16#29f7# => X"18400001",
		16#29f8# => X"a8428768",
		16#29f9# => X"03ffffe4",
		16#29fa# => X"85620000",
		16#29fb# => X"d7e117f4",
		16#29fc# => X"9c800000",
		16#29fd# => X"d7e14ffc",
		16#29fe# => X"d7e177f8",
		16#29ff# => X"9c21ffe4",
		16#2a00# => X"a8430000",
		16#2a01# => X"e4232000",
		16#2a02# => X"0c000018",
		16#2a03# => X"d4012004",
		16#2a04# => X"9c800003",
		16#2a05# => X"9dc0001e",
		16#2a06# => X"d4012000",
		16#2a07# => X"d4017008",
		16#2a08# => X"04000734",
		16#2a09# => X"d401180c",
		16#2a0a# => X"9d6bffff",
		16#2a0b# => X"bd6b0000",
		16#2a0c# => X"0c000017",
		16#2a0d# => X"bc0b0000",
		16#2a0e# => X"10000005",
		16#2a0f# => X"e0425808",
		16#2a10# => X"e16e5802",
		16#2a11# => X"d401100c",
		16#2a12# => X"d4015808",
		16#2a13# => X"07fffccd",
		16#2a14# => X"a8610000",
		16#2a15# => X"9c21001c",
		16#2a16# => X"8521fffc",
		16#2a17# => X"8441fff4",
		16#2a18# => X"44004800",
		16#2a19# => X"85c1fff8",
		16#2a1a# => X"9c400002",
		16#2a1b# => X"a8610000",
		16#2a1c# => X"07fffcc4",
		16#2a1d# => X"d4011000",
		16#2a1e# => X"9c21001c",
		16#2a1f# => X"8521fffc",
		16#2a20# => X"8441fff4",
		16#2a21# => X"44004800",
		16#2a22# => X"85c1fff8",
		16#2a23# => X"e0605802",
		16#2a24# => X"9ca00001",
		16#2a25# => X"e0821848",
		16#2a26# => X"e0651808",
		16#2a27# => X"e16e5802",
		16#2a28# => X"9c63ffff",
		16#2a29# => X"d4015808",
		16#2a2a# => X"e0431003",
		16#2a2b# => X"e0601002",
		16#2a2c# => X"e0431004",
		16#2a2d# => X"a8610000",
		16#2a2e# => X"b842005f",
		16#2a2f# => X"e0422004",
		16#2a30# => X"07fffcb0",
		16#2a31# => X"d401100c",
		16#2a32# => X"9c21001c",
		16#2a33# => X"8521fffc",
		16#2a34# => X"8441fff4",
		16#2a35# => X"44004800",
		16#2a36# => X"85c1fff8",
		16#2a37# => X"d7e14ffc",
		16#2a38# => X"9c21ffe8",
		16#2a39# => X"d4011810",
		16#2a3a# => X"a8810000",
		16#2a3b# => X"07fffd12",
		16#2a3c# => X"9c610010",
		16#2a3d# => X"84610000",
		16#2a3e# => X"bc030002",
		16#2a3f# => X"10000012",
		16#2a40# => X"9d600000",
		16#2a41# => X"bca30001",
		16#2a42# => X"1000000f",
		16#2a43# => X"bc230004",
		16#2a44# => X"0c00001d",
		16#2a45# => X"84610008",
		16#2a46# => X"bd830000",
		16#2a47# => X"1000000a",
		16#2a48# => X"bda3001e",
		16#2a49# => X"1000000c",
		16#2a4a# => X"15000000",
		16#2a4b# => X"84610004",
		16#2a4c# => X"bc030000",
		16#2a4d# => X"0c000018",
		16#2a4e# => X"15000000",
		16#2a4f# => X"19607fff",
		16#2a50# => X"a96bffff",
		16#2a51# => X"9c210018",
		16#2a52# => X"8521fffc",
		16#2a53# => X"44004800",
		16#2a54# => X"15000000",
		16#2a55# => X"9d60001e",
		16#2a56# => X"e06b1802",
		16#2a57# => X"8561000c",
		16#2a58# => X"e16b1848",
		16#2a59# => X"84610004",
		16#2a5a# => X"bc030000",
		16#2a5b# => X"13fffff6",
		16#2a5c# => X"15000000",
		16#2a5d# => X"9c210018",
		16#2a5e# => X"8521fffc",
		16#2a5f# => X"44004800",
		16#2a60# => X"e1605802",
		16#2a61# => X"84610004",
		16#2a62# => X"e4035800",
		16#2a63# => X"13ffffec",
		16#2a64# => X"15000000",
		16#2a65# => X"9c210018",
		16#2a66# => X"8521fffc",
		16#2a67# => X"44004800",
		16#2a68# => X"19608000",
		16#2a69# => X"d7e14ffc",
		16#2a6a# => X"d7e117f8",
		16#2a6b# => X"9c21ffe4",
		16#2a6c# => X"d4011810",
		16#2a6d# => X"a8810000",
		16#2a6e# => X"07fffcdf",
		16#2a6f# => X"9c610010",
		16#2a70# => X"84810004",
		16#2a71# => X"a8610000",
		16#2a72# => X"e0402002",
		16#2a73# => X"e0422004",
		16#2a74# => X"ac42ffff",
		16#2a75# => X"b842005f",
		16#2a76# => X"07fffc6a",
		16#2a77# => X"d4011004",
		16#2a78# => X"9c21001c",
		16#2a79# => X"8521fffc",
		16#2a7a# => X"44004800",
		16#2a7b# => X"8441fff8",
		16#2a7c# => X"d7e14ffc",
		16#2a7d# => X"9c21ffec",
		16#2a7e# => X"d4011800",
		16#2a7f# => X"a8610000",
		16#2a80# => X"d4012004",
		16#2a81# => X"d4012808",
		16#2a82# => X"07fffc5e",
		16#2a83# => X"d401300c",
		16#2a84# => X"9c210014",
		16#2a85# => X"8521fffc",
		16#2a86# => X"44004800",
		16#2a87# => X"15000000",
		16#2a88# => X"d7e14ffc",
		16#2a89# => X"d7e117f8",
		16#2a8a# => X"9c21ffe4",
		16#2a8b# => X"d4011810",
		16#2a8c# => X"a8810000",
		16#2a8d# => X"07fffcc0",
		16#2a8e# => X"9c610010",
		16#2a8f# => X"84e1000c",
		16#2a90# => X"84610000",
		16#2a91# => X"b8c70042",
		16#2a92# => X"b8e7001e",
		16#2a93# => X"84810004",
		16#2a94# => X"04000636",
		16#2a95# => X"84a10008",
		16#2a96# => X"9c21001c",
		16#2a97# => X"a84b0000",
		16#2a98# => X"a86c0000",
		16#2a99# => X"8521fffc",
		16#2a9a# => X"e1620004",
		16#2a9b# => X"e1830004",
		16#2a9c# => X"44004800",
		16#2a9d# => X"8441fff8",
		16#2a9e# => X"d7e117f8",
		16#2a9f# => X"d7e177fc",
		16#2aa0# => X"84430000",
		16#2aa1# => X"9c21fff8",
		16#2aa2# => X"bca20001",
		16#2aa3# => X"1000008c",
		16#2aa4# => X"a9630000",
		16#2aa5# => X"84640000",
		16#2aa6# => X"bca30001",
		16#2aa7# => X"100000cf",
		16#2aa8# => X"bc220004",
		16#2aa9# => X"0c000109",
		16#2aaa# => X"bc030004",
		16#2aab# => X"100000cb",
		16#2aac# => X"bc230002",
		16#2aad# => X"0c00009a",
		16#2aae# => X"bc020002",
		16#2aaf# => X"100000c7",
		16#2ab0# => X"15000000",
		16#2ab1# => X"858b0008",
		16#2ab2# => X"85e40008",
		16#2ab3# => X"84cb000c",
		16#2ab4# => X"84eb0010",
		16#2ab5# => X"e1ac7802",
		16#2ab6# => X"8444000c",
		16#2ab7# => X"84640010",
		16#2ab8# => X"ba2d009f",
		16#2ab9# => X"e1116805",
		16#2aba# => X"e1088802",
		16#2abb# => X"bd48003f",
		16#2abc# => X"10000077",
		16#2abd# => X"e5ac7800",
		16#2abe# => X"bdad0000",
		16#2abf# => X"100000bc",
		16#2ac0# => X"bc0d0000",
		16#2ac1# => X"9da8ffe0",
		16#2ac2# => X"bd8d0000",
		16#2ac3# => X"100000d4",
		16#2ac4# => X"a9c20000",
		16#2ac5# => X"9ea00000",
		16#2ac6# => X"e1ee6848",
		16#2ac7# => X"bd8d0000",
		16#2ac8# => X"100000dc",
		16#2ac9# => X"9e200001",
		16#2aca# => X"9d000000",
		16#2acb# => X"e1b16808",
		16#2acc# => X"9e28ffff",
		16#2acd# => X"e4914000",
		16#2ace# => X"10000003",
		16#2acf# => X"9e600001",
		16#2ad0# => X"9e600000",
		16#2ad1# => X"9d0dffff",
		16#2ad2# => X"e2311803",
		16#2ad3# => X"e1134000",
		16#2ad4# => X"e1081003",
		16#2ad5# => X"a8550000",
		16#2ad6# => X"e1088804",
		16#2ad7# => X"e1a04002",
		16#2ad8# => X"e10d4004",
		16#2ad9# => X"b908005f",
		16#2ada# => X"e1e87804",
		16#2adb# => X"a86f0000",
		16#2adc# => X"850b0004",
		16#2add# => X"84840004",
		16#2ade# => X"e4082000",
		16#2adf# => X"1000005d",
		16#2ae0# => X"e0833800",
		16#2ae1# => X"bc080000",
		16#2ae2# => X"1000007f",
		16#2ae3# => X"e0871802",
		16#2ae4# => X"e0833802",
		16#2ae5# => X"e4441800",
		16#2ae6# => X"10000003",
		16#2ae7# => X"9d000001",
		16#2ae8# => X"9d000000",
		16#2ae9# => X"e0623002",
		16#2aea# => X"e0634002",
		16#2aeb# => X"bd830000",
		16#2aec# => X"1000007f",
		16#2aed# => X"9c400001",
		16#2aee# => X"9d600000",
		16#2aef# => X"d4056008",
		16#2af0# => X"d4055804",
		16#2af1# => X"d405180c",
		16#2af2# => X"d4052010",
		16#2af3# => X"9cc4ffff",
		16#2af4# => X"e4862000",
		16#2af5# => X"10000003",
		16#2af6# => X"9c400001",
		16#2af7# => X"9c400000",
		16#2af8# => X"9ce3ffff",
		16#2af9# => X"19a00fff",
		16#2afa# => X"e0423800",
		16#2afb# => X"a9adffff",
		16#2afc# => X"e4426800",
		16#2afd# => X"10000020",
		16#2afe# => X"e4226800",
		16#2aff# => X"0c0000a1",
		16#2b00# => X"bc46fffe",
		16#2b01# => X"00000004",
		16#2b02# => X"84450008",
		16#2b03# => X"0c00005a",
		16#2b04# => X"bc4bfffe",
		16#2b05# => X"e0c42000",
		16#2b06# => X"e0631800",
		16#2b07# => X"9d66ffff",
		16#2b08# => X"e4862000",
		16#2b09# => X"10000003",
		16#2b0a# => X"9d000001",
		16#2b0b# => X"9d000000",
		16#2b0c# => X"e0681800",
		16#2b0d# => X"9ce00001",
		16#2b0e# => X"e48b3000",
		16#2b0f# => X"9d03ffff",
		16#2b10# => X"a8860000",
		16#2b11# => X"10000003",
		16#2b12# => X"9c42ffff",
		16#2b13# => X"9ce00000",
		16#2b14# => X"e0e74000",
		16#2b15# => X"19000fff",
		16#2b16# => X"a908ffff",
		16#2b17# => X"e4474000",
		16#2b18# => X"0fffffeb",
		16#2b19# => X"e4274000",
		16#2b1a# => X"d405180c",
		16#2b1b# => X"d4053010",
		16#2b1c# => X"d4051008",
		16#2b1d# => X"19a01fff",
		16#2b1e# => X"9c400003",
		16#2b1f# => X"a9adffff",
		16#2b20# => X"e4436800",
		16#2b21# => X"0c00000d",
		16#2b22# => X"d4051000",
		16#2b23# => X"b8e3001f",
		16#2b24# => X"b8440041",
		16#2b25# => X"84c50008",
		16#2b26# => X"a4840001",
		16#2b27# => X"e0471004",
		16#2b28# => X"b8630041",
		16#2b29# => X"e0441004",
		16#2b2a# => X"9cc60001",
		16#2b2b# => X"d405180c",
		16#2b2c# => X"d4051010",
		16#2b2d# => X"d4053008",
		16#2b2e# => X"a9650000",
		16#2b2f# => X"9c210008",
		16#2b30# => X"8441fff8",
		16#2b31# => X"44004800",
		16#2b32# => X"85c1fffc",
		16#2b33# => X"10000026",
		16#2b34# => X"15000000",
		16#2b35# => X"850b0004",
		16#2b36# => X"84840004",
		16#2b37# => X"9c400000",
		16#2b38# => X"e4082000",
		16#2b39# => X"0fffffa8",
		16#2b3a# => X"9c600000",
		16#2b3b# => X"e0833800",
		16#2b3c# => X"d4054004",
		16#2b3d# => X"d4056008",
		16#2b3e# => X"e4841800",
		16#2b3f# => X"10000003",
		16#2b40# => X"9d000001",
		16#2b41# => X"9d000000",
		16#2b42# => X"e0423000",
		16#2b43# => X"d4052010",
		16#2b44# => X"e0681000",
		16#2b45# => X"03ffffd8",
		16#2b46# => X"d405180c",
		16#2b47# => X"bc220002",
		16#2b48# => X"13ffffe7",
		16#2b49# => X"15000000",
		16#2b4a# => X"d4051000",
		16#2b4b# => X"844b0004",
		16#2b4c# => X"d4051004",
		16#2b4d# => X"844b0008",
		16#2b4e# => X"d4051008",
		16#2b4f# => X"844b000c",
		16#2b50# => X"d405100c",
		16#2b51# => X"844b0010",
		16#2b52# => X"d4051010",
		16#2b53# => X"844b0004",
		16#2b54# => X"84640004",
		16#2b55# => X"a9650000",
		16#2b56# => X"e0431003",
		16#2b57# => X"03ffffd8",
		16#2b58# => X"d4051004",
		16#2b59# => X"a98f0000",
		16#2b5a# => X"9cc00000",
		16#2b5b# => X"03ffff81",
		16#2b5c# => X"9ce00000",
		16#2b5d# => X"0fffffa8",
		16#2b5e# => X"15000000",
		16#2b5f# => X"03ffffbc",
		16#2b60# => X"d405180c",
		16#2b61# => X"e4443800",
		16#2b62# => X"10000003",
		16#2b63# => X"9d600001",
		16#2b64# => X"a9680000",
		16#2b65# => X"e0661002",
		16#2b66# => X"e0635802",
		16#2b67# => X"bd830000",
		16#2b68# => X"0fffff87",
		16#2b69# => X"9d600000",
		16#2b6a# => X"9c400001",
		16#2b6b# => X"e0802002",
		16#2b6c# => X"d4051004",
		16#2b6d# => X"bc440000",
		16#2b6e# => X"10000003",
		16#2b6f# => X"d4056008",
		16#2b70# => X"9c400000",
		16#2b71# => X"e0601802",
		16#2b72# => X"d4052010",
		16#2b73# => X"e0631002",
		16#2b74# => X"03ffff7f",
		16#2b75# => X"d405180c",
		16#2b76# => X"9c210008",
		16#2b77# => X"a9640000",
		16#2b78# => X"8441fff8",
		16#2b79# => X"44004800",
		16#2b7a# => X"85c1fffc",
		16#2b7b# => X"13ffff61",
		16#2b7c# => X"9da8ffe0",
		16#2b7d# => X"bd8d0000",
		16#2b7e# => X"1000002c",
		16#2b7f# => X"e18c4000",
		16#2b80# => X"e1e66848",
		16#2b81# => X"9ea00000",
		16#2b82# => X"bd8d0000",
		16#2b83# => X"10000024",
		16#2b84# => X"9e200001",
		16#2b85# => X"9d000000",
		16#2b86# => X"e1b16808",
		16#2b87# => X"9e28ffff",
		16#2b88# => X"e4914000",
		16#2b89# => X"10000003",
		16#2b8a# => X"9e600001",
		16#2b8b# => X"9e600000",
		16#2b8c# => X"9d0dffff",
		16#2b8d# => X"e2313803",
		16#2b8e# => X"e1134000",
		16#2b8f# => X"e1083003",
		16#2b90# => X"a8d50000",
		16#2b91# => X"e1088804",
		16#2b92# => X"e1a04002",
		16#2b93# => X"e10d4004",
		16#2b94# => X"b908005f",
		16#2b95# => X"03ffff47",
		16#2b96# => X"e0e87804",
		16#2b97# => X"9e20001f",
		16#2b98# => X"ba6e0001",
		16#2b99# => X"e2314002",
		16#2b9a# => X"e1e34048",
		16#2b9b# => X"e2338808",
		16#2b9c# => X"a9c20000",
		16#2b9d# => X"e1f17804",
		16#2b9e# => X"03ffff29",
		16#2b9f# => X"e2ae4048",
		16#2ba0# => X"0fffff61",
		16#2ba1# => X"15000000",
		16#2ba2# => X"03ffff7c",
		16#2ba3# => X"19a01fff",
		16#2ba4# => X"9da00000",
		16#2ba5# => X"03ffff27",
		16#2ba6# => X"e1114008",
		16#2ba7# => X"9da00000",
		16#2ba8# => X"03ffffdf",
		16#2ba9# => X"e1114008",
		16#2baa# => X"9e20001f",
		16#2bab# => X"ba660001",
		16#2bac# => X"e2314002",
		16#2bad# => X"e1e74048",
		16#2bae# => X"e2338808",
		16#2baf# => X"e2a64048",
		16#2bb0# => X"03ffffd2",
		16#2bb1# => X"e1f17804",
		16#2bb2# => X"bc230004",
		16#2bb3# => X"13ffff7c",
		16#2bb4# => X"15000000",
		16#2bb5# => X"846b0004",
		16#2bb6# => X"84440004",
		16#2bb7# => X"e4231000",
		16#2bb8# => X"0fffff77",
		16#2bb9# => X"15000000",
		16#2bba# => X"19600001",
		16#2bbb# => X"03ffff74",
		16#2bbc# => X"a96b877c",
		16#2bbd# => X"d7e187ec",
		16#2bbe# => X"d7e14ffc",
		16#2bbf# => X"d7e117e4",
		16#2bc0# => X"d7e177e8",
		16#2bc1# => X"d7e197f0",
		16#2bc2# => X"d7e1a7f4",
		16#2bc3# => X"d7e1b7f8",
		16#2bc4# => X"84830000",
		16#2bc5# => X"9c21ffdc",
		16#2bc6# => X"8443000c",
		16#2bc7# => X"85c30010",
		16#2bc8# => X"bc440001",
		16#2bc9# => X"0c000051",
		16#2bca# => X"86030004",
		16#2bcb# => X"bc040004",
		16#2bcc# => X"10000049",
		16#2bcd# => X"bc040002",
		16#2bce# => X"1000002a",
		16#2bcf# => X"e0827004",
		16#2bd0# => X"bc040000",
		16#2bd1# => X"10000027",
		16#2bd2# => X"15000000",
		16#2bd3# => X"84630008",
		16#2bd4# => X"bd63fc02",
		16#2bd5# => X"0c00004e",
		16#2bd6# => X"bd4303ff",
		16#2bd7# => X"1000003e",
		16#2bd8# => X"a48e00ff",
		16#2bd9# => X"bc240080",
		16#2bda# => X"0c000031",
		16#2bdb# => X"9c6303ff",
		16#2bdc# => X"9c8e007f",
		16#2bdd# => X"e4847000",
		16#2bde# => X"0c000035",
		16#2bdf# => X"9ca00001",
		16#2be0# => X"e0451000",
		16#2be1# => X"a9c40000",
		16#2be2# => X"18a01fff",
		16#2be3# => X"a8a5ffff",
		16#2be4# => X"e4422800",
		16#2be5# => X"0c000006",
		16#2be6# => X"b882001f",
		16#2be7# => X"b9ce0041",
		16#2be8# => X"b8420041",
		16#2be9# => X"9c630001",
		16#2bea# => X"e1c47004",
		16#2beb# => X"a4a307ff",
		16#2bec# => X"1900000f",
		16#2bed# => X"b8e20048",
		16#2bee# => X"b8a50014",
		16#2bef# => X"a908ffff",
		16#2bf0# => X"b8820018",
		16#2bf1# => X"b9ce0048",
		16#2bf2# => X"a8450000",
		16#2bf3# => X"e0a74003",
		16#2bf4# => X"9ce00000",
		16#2bf5# => X"e0c47004",
		16#2bf6# => X"00000006",
		16#2bf7# => X"a8670000",
		16#2bf8# => X"9c400000",
		16#2bf9# => X"9c600000",
		16#2bfa# => X"e0a20004",
		16#2bfb# => X"e0c30004",
		16#2bfc# => X"b890001f",
		16#2bfd# => X"9c210024",
		16#2bfe# => X"e0e51004",
		16#2bff# => X"8521fffc",
		16#2c00# => X"e0461804",
		16#2c01# => X"e0672004",
		16#2c02# => X"a9820000",
		16#2c03# => X"a9630000",
		16#2c04# => X"8441ffe4",
		16#2c05# => X"85c1ffe8",
		16#2c06# => X"8601ffec",
		16#2c07# => X"8641fff0",
		16#2c08# => X"8681fff4",
		16#2c09# => X"44004800",
		16#2c0a# => X"86c1fff8",
		16#2c0b# => X"a48e0100",
		16#2c0c# => X"bc040000",
		16#2c0d# => X"13ffffd6",
		16#2c0e# => X"18a01fff",
		16#2c0f# => X"9c8e0080",
		16#2c10# => X"e4847000",
		16#2c11# => X"13ffffcf",
		16#2c12# => X"9ca00001",
		16#2c13# => X"03ffffcd",
		16#2c14# => X"9ca00000",
		16#2c15# => X"18407ff0",
		16#2c16# => X"9c600000",
		16#2c17# => X"9ca00000",
		16#2c18# => X"03ffffe4",
		16#2c19# => X"9cc00000",
		16#2c1a# => X"18600008",
		16#2c1b# => X"1880000f",
		16#2c1c# => X"e0421804",
		16#2c1d# => X"a884ffff",
		16#2c1e# => X"9c600000",
		16#2c1f# => X"e0a22003",
		16#2c20# => X"a8ce0000",
		16#2c21# => X"03ffffdb",
		16#2c22# => X"18407ff0",
		16#2c23# => X"9e40fc02",
		16#2c24# => X"9ce00000",
		16#2c25# => X"9d000000",
		16#2c26# => X"e2521802",
		16#2c27# => X"d4013800",
		16#2c28# => X"d4014004",
		16#2c29# => X"bd520038",
		16#2c2a# => X"10000046",
		16#2c2b# => X"85010004",
		16#2c2c# => X"a8620000",
		16#2c2d# => X"a88e0000",
		16#2c2e# => X"040004e6",
		16#2c2f# => X"a8b20000",
		16#2c30# => X"a8b20000",
		16#2c31# => X"9c600000",
		16#2c32# => X"9c800001",
		16#2c33# => X"aacb0000",
		16#2c34# => X"040004f4",
		16#2c35# => X"aa8c0000",
		16#2c36# => X"9c800001",
		16#2c37# => X"a86b0000",
		16#2c38# => X"bc2c0000",
		16#2c39# => X"10000003",
		16#2c3a# => X"9cacffff",
		16#2c3b# => X"9c800000",
		16#2c3c# => X"9c63ffff",
		16#2c3d# => X"e1c57003",
		16#2c3e# => X"e0841800",
		16#2c3f# => X"d401b000",
		16#2c40# => X"e0441003",
		16#2c41# => X"e0427004",
		16#2c42# => X"e0601002",
		16#2c43# => X"e0431004",
		16#2c44# => X"b842005f",
		16#2c45# => X"e282a004",
		16#2c46# => X"a45400ff",
		16#2c47# => X"bc220080",
		16#2c48# => X"10000027",
		16#2c49# => X"d401a004",
		16#2c4a# => X"a4540100",
		16#2c4b# => X"bc020000",
		16#2c4c# => X"1000000e",
		16#2c4d# => X"85010000",
		16#2c4e# => X"9c540080",
		16#2c4f# => X"e482a000",
		16#2c50# => X"0c000024",
		16#2c51# => X"9c600001",
		16#2c52# => X"84e10000",
		16#2c53# => X"a8820000",
		16#2c54# => X"e0a33800",
		16#2c55# => X"a8640000",
		16#2c56# => X"a8450000",
		16#2c57# => X"d4011000",
		16#2c58# => X"d4011804",
		16#2c59# => X"85010000",
		16#2c5a# => X"84a10004",
		16#2c5b# => X"b8e80018",
		16#2c5c# => X"b8850048",
		16#2c5d# => X"b8480048",
		16#2c5e# => X"1900000f",
		16#2c5f# => X"e0c72004",
		16#2c60# => X"18e00fff",
		16#2c61# => X"a908ffff",
		16#2c62# => X"84810000",
		16#2c63# => X"a8e7ffff",
		16#2c64# => X"e0a24003",
		16#2c65# => X"e4443800",
		16#2c66# => X"10000003",
		16#2c67# => X"9c600001",
		16#2c68# => X"9c600000",
		16#2c69# => X"a48307ff",
		16#2c6a# => X"b8840014",
		16#2c6b# => X"a8440000",
		16#2c6c# => X"9c800000",
		16#2c6d# => X"03ffff8f",
		16#2c6e# => X"a8640000",
		16#2c6f# => X"85010004",
		16#2c70# => X"9c48007f",
		16#2c71# => X"e4824000",
		16#2c72# => X"13ffffe0",
		16#2c73# => X"9c600001",
		16#2c74# => X"03ffffde",
		16#2c75# => X"9c600000",
		16#2c76# => X"d7e117fc",
		16#2c77# => X"1840000f",
		16#2c78# => X"84c30000",
		16#2c79# => X"84a30004",
		16#2c7a# => X"b8e60054",
		16#2c7b# => X"b906005f",
		16#2c7c# => X"a842ffff",
		16#2c7d# => X"a4e707ff",
		16#2c7e# => X"d4044004",
		16#2c7f# => X"9c21fffc",
		16#2c80# => X"bc270000",
		16#2c81# => X"10000022",
		16#2c82# => X"e0661003",
		16#2c83# => X"e0c32804",
		16#2c84# => X"bc260000",
		16#2c85# => X"0c00002f",
		16#2c86# => X"b8c50058",
		16#2c87# => X"b8630008",
		16#2c88# => X"9ce0fc02",
		16#2c89# => X"b8a50008",
		16#2c8a# => X"e0661804",
		16#2c8b# => X"9cc00003",
		16#2c8c# => X"d4043808",
		16#2c8d# => X"d4043000",
		16#2c8e# => X"9cc0fc01",
		16#2c8f# => X"e0e52800",
		16#2c90# => X"e0631800",
		16#2c91# => X"e4872800",
		16#2c92# => X"10000003",
		16#2c93# => X"9d000001",
		16#2c94# => X"9d000000",
		16#2c95# => X"18400fff",
		16#2c96# => X"e0681800",
		16#2c97# => X"a842ffff",
		16#2c98# => X"a9660000",
		16#2c99# => X"a8a70000",
		16#2c9a# => X"e4431000",
		16#2c9b# => X"0ffffff4",
		16#2c9c# => X"9cc6ffff",
		16#2c9d# => X"9c210004",
		16#2c9e# => X"d4045808",
		16#2c9f# => X"d404180c",
		16#2ca0# => X"d4043810",
		16#2ca1# => X"44004800",
		16#2ca2# => X"8441fffc",
		16#2ca3# => X"bc2707ff",
		16#2ca4# => X"0c000015",
		16#2ca5# => X"9ce7fc01",
		16#2ca6# => X"b8c50058",
		16#2ca7# => X"b8630008",
		16#2ca8# => X"18401000",
		16#2ca9# => X"e0661804",
		16#2caa# => X"b8a50008",
		16#2cab# => X"e0631004",
		16#2cac# => X"d4043808",
		16#2cad# => X"9cc00003",
		16#2cae# => X"d4043000",
		16#2caf# => X"d404180c",
		16#2cb0# => X"d4042810",
		16#2cb1# => X"9c210004",
		16#2cb2# => X"44004800",
		16#2cb3# => X"8441fffc",
		16#2cb4# => X"9c600002",
		16#2cb5# => X"9c210004",
		16#2cb6# => X"d4041800",
		16#2cb7# => X"44004800",
		16#2cb8# => X"8441fffc",
		16#2cb9# => X"e0e32804",
		16#2cba# => X"bc270000",
		16#2cbb# => X"0c00000a",
		16#2cbc# => X"15000000",
		16#2cbd# => X"18400008",
		16#2cbe# => X"e0c61003",
		16#2cbf# => X"bc060000",
		16#2cc0# => X"13ffffee",
		16#2cc1# => X"15000000",
		16#2cc2# => X"9cc00001",
		16#2cc3# => X"03ffffec",
		16#2cc4# => X"d4043000",
		16#2cc5# => X"9c600004",
		16#2cc6# => X"03ffffeb",
		16#2cc7# => X"d4041800",
		16#2cc8# => X"d7e14ffc",
		16#2cc9# => X"d7e117f4",
		16#2cca# => X"d7e177f8",
		16#2ccb# => X"9c21ffa8",
		16#2ccc# => X"9dc10028",
		16#2ccd# => X"d4011844",
		16#2cce# => X"d4012048",
		16#2ccf# => X"9c610044",
		16#2cd0# => X"a88e0000",
		16#2cd1# => X"d401283c",
		16#2cd2# => X"d4013040",
		16#2cd3# => X"07ffffa3",
		16#2cd4# => X"9c410014",
		16#2cd5# => X"9c61003c",
		16#2cd6# => X"07ffffa0",
		16#2cd7# => X"a8820000",
		16#2cd8# => X"a86e0000",
		16#2cd9# => X"a8820000",
		16#2cda# => X"07fffdc4",
		16#2cdb# => X"a8a10000",
		16#2cdc# => X"07fffee1",
		16#2cdd# => X"a86b0000",
		16#2cde# => X"9c210058",
		16#2cdf# => X"a84b0000",
		16#2ce0# => X"a86c0000",
		16#2ce1# => X"8521fffc",
		16#2ce2# => X"e1620004",
		16#2ce3# => X"e1830004",
		16#2ce4# => X"85c1fff8",
		16#2ce5# => X"44004800",
		16#2ce6# => X"8441fff4",
		16#2ce7# => X"d7e14ffc",
		16#2ce8# => X"d7e117f4",
		16#2ce9# => X"d7e177f8",
		16#2cea# => X"9c21ffa8",
		16#2ceb# => X"9c410028",
		16#2cec# => X"d4011844",
		16#2ced# => X"d4012048",
		16#2cee# => X"9c610044",
		16#2cef# => X"a8820000",
		16#2cf0# => X"d401283c",
		16#2cf1# => X"d4013040",
		16#2cf2# => X"07ffff84",
		16#2cf3# => X"9dc10014",
		16#2cf4# => X"9c61003c",
		16#2cf5# => X"07ffff81",
		16#2cf6# => X"a88e0000",
		16#2cf7# => X"84c10018",
		16#2cf8# => X"a88e0000",
		16#2cf9# => X"acc60001",
		16#2cfa# => X"a8a10000",
		16#2cfb# => X"a8620000",
		16#2cfc# => X"07fffda2",
		16#2cfd# => X"d4013018",
		16#2cfe# => X"07fffebf",
		16#2cff# => X"a86b0000",
		16#2d00# => X"9c210058",
		16#2d01# => X"a84b0000",
		16#2d02# => X"a86c0000",
		16#2d03# => X"8521fffc",
		16#2d04# => X"e1620004",
		16#2d05# => X"e1830004",
		16#2d06# => X"85c1fff8",
		16#2d07# => X"44004800",
		16#2d08# => X"8441fff4",
		16#2d09# => X"d7e14ffc",
		16#2d0a# => X"d7e117dc",
		16#2d0b# => X"d7e177e0",
		16#2d0c# => X"d7e187e4",
		16#2d0d# => X"d7e197e8",
		16#2d0e# => X"d7e1a7ec",
		16#2d0f# => X"d7e1b7f0",
		16#2d10# => X"d7e1c7f4",
		16#2d11# => X"d7e1d7f8",
		16#2d12# => X"9c21ff90",
		16#2d13# => X"9dc10028",
		16#2d14# => X"d4011844",
		16#2d15# => X"d4012048",
		16#2d16# => X"9c610044",
		16#2d17# => X"a88e0000",
		16#2d18# => X"d401283c",
		16#2d19# => X"d4013040",
		16#2d1a# => X"07ffff5c",
		16#2d1b# => X"9e010014",
		16#2d1c# => X"9c61003c",
		16#2d1d# => X"07ffff59",
		16#2d1e# => X"a8900000",
		16#2d1f# => X"84410028",
		16#2d20# => X"bc420001",
		16#2d21# => X"0c0000c7",
		16#2d22# => X"84a10014",
		16#2d23# => X"bc450001",
		16#2d24# => X"0c0000df",
		16#2d25# => X"bc220004",
		16#2d26# => X"0c0000be",
		16#2d27# => X"bc250004",
		16#2d28# => X"0c0000d7",
		16#2d29# => X"bc220002",
		16#2d2a# => X"0c0000be",
		16#2d2b# => X"bc250002",
		16#2d2c# => X"0c0000d7",
		16#2d2d# => X"84410038",
		16#2d2e# => X"9c600000",
		16#2d2f# => X"86010024",
		16#2d30# => X"a8a30000",
		16#2d31# => X"a8820000",
		16#2d32# => X"a8d00000",
		16#2d33# => X"040003c4",
		16#2d34# => X"86810020",
		16#2d35# => X"9c600000",
		16#2d36# => X"a8940000",
		16#2d37# => X"a8a30000",
		16#2d38# => X"a8c20000",
		16#2d39# => X"a9cb0000",
		16#2d3a# => X"040003bd",
		16#2d3b# => X"ab0c0000",
		16#2d3c# => X"9c600000",
		16#2d3d# => X"87410034",
		16#2d3e# => X"a8a30000",
		16#2d3f# => X"a8d40000",
		16#2d40# => X"a89a0000",
		16#2d41# => X"aa4c0000",
		16#2d42# => X"040003b5",
		16#2d43# => X"a84b0000",
		16#2d44# => X"9c600000",
		16#2d45# => X"a89a0000",
		16#2d46# => X"a8a30000",
		16#2d47# => X"a8d00000",
		16#2d48# => X"aa8b0000",
		16#2d49# => X"040003ae",
		16#2d4a# => X"aacc0000",
		16#2d4b# => X"e0ac9000",
		16#2d4c# => X"a90b0000",
		16#2d4d# => X"e4856000",
		16#2d4e# => X"0c00006d",
		16#2d4f# => X"9da00001",
		16#2d50# => X"e0e81000",
		16#2d51# => X"e0ed3800",
		16#2d52# => X"e4423800",
		16#2d53# => X"0c000063",
		16#2d54# => X"e4223800",
		16#2d55# => X"9c400001",
		16#2d56# => X"9c600000",
		16#2d57# => X"e0a57000",
		16#2d58# => X"e44e2800",
		16#2d59# => X"0c000009",
		16#2d5a# => X"a8d80000",
		16#2d5b# => X"9c830001",
		16#2d5c# => X"e4841800",
		16#2d5d# => X"0c000081",
		16#2d5e# => X"9d000001",
		16#2d5f# => X"e1081000",
		16#2d60# => X"a8640000",
		16#2d61# => X"a8480000",
		16#2d62# => X"e187b000",
		16#2d63# => X"e48c3800",
		16#2d64# => X"10000003",
		16#2d65# => X"9c800001",
		16#2d66# => X"9c800000",
		16#2d67# => X"e10c1800",
		16#2d68# => X"e084a000",
		16#2d69# => X"e4886000",
		16#2d6a# => X"10000003",
		16#2d6b# => X"9da00001",
		16#2d6c# => X"9da00000",
		16#2d6d# => X"84e10018",
		16#2d6e# => X"8581002c",
		16#2d6f# => X"85c1001c",
		16#2d70# => X"e18c3805",
		16#2d71# => X"84e10030",
		16#2d72# => X"e1606002",
		16#2d73# => X"e0ee3800",
		16#2d74# => X"e18b6004",
		16#2d75# => X"e0841000",
		16#2d76# => X"b98c005f",
		16#2d77# => X"9c670004",
		16#2d78# => X"18401fff",
		16#2d79# => X"e08d2000",
		16#2d7a# => X"d4011808",
		16#2d7b# => X"a842ffff",
		16#2d7c# => X"d4016004",
		16#2d7d# => X"e4441000",
		16#2d7e# => X"0c000017",
		16#2d7f# => X"a8680000",
		16#2d80# => X"9ce70005",
		16#2d81# => X"b9030041",
		16#2d82# => X"a4630001",
		16#2d83# => X"b964001f",
		16#2d84# => X"b985001f",
		16#2d85# => X"b8460041",
		16#2d86# => X"b9a50041",
		16#2d87# => X"b8840041",
		16#2d88# => X"bc030000",
		16#2d89# => X"10000005",
		16#2d8a# => X"a9e70000",
		16#2d8b# => X"18608000",
		16#2d8c# => X"e0cc1004",
		16#2d8d# => X"e0ad1804",
		16#2d8e# => X"e06b4004",
		16#2d8f# => X"19001fff",
		16#2d90# => X"a908ffff",
		16#2d91# => X"e4444000",
		16#2d92# => X"13ffffef",
		16#2d93# => X"9ce70001",
		16#2d94# => X"d4017808",
		16#2d95# => X"19600fff",
		16#2d96# => X"a96bffff",
		16#2d97# => X"e4445800",
		16#2d98# => X"1000002c",
		16#2d99# => X"84e10008",
		16#2d9a# => X"0000000d",
		16#2d9b# => X"e1631800",
		16#2d9c# => X"e4883000",
		16#2d9d# => X"10000003",
		16#2d9e# => X"9ca00001",
		16#2d9f# => X"9ca00000",
		16#2da0# => X"18400fff",
		16#2da1# => X"a8c80000",
		16#2da2# => X"a842ffff",
		16#2da3# => X"e44b1000",
		16#2da4# => X"1000001f",
		16#2da5# => X"e0a56800",
		16#2da6# => X"e1631800",
		16#2da7# => X"e0842000",
		16#2da8# => X"e1063000",
		16#2da9# => X"e1a52800",
		16#2daa# => X"9d800001",
		16#2dab# => X"e48b1800",
		16#2dac# => X"10000003",
		16#2dad# => X"9ce7ffff",
		16#2dae# => X"9d800000",
		16#2daf# => X"e08c2000",
		16#2db0# => X"a86b0000",
		16#2db1# => X"bd850000",
		16#2db2# => X"0fffffea",
		16#2db3# => X"a9640000",
		16#2db4# => X"03ffffe8",
		16#2db5# => X"a8630001",
		16#2db6# => X"0c00002a",
		16#2db7# => X"e4522800",
		16#2db8# => X"9c400000",
		16#2db9# => X"03ffff9e",
		16#2dba# => X"9c600000",
		16#2dbb# => X"9da00000",
		16#2dbc# => X"e0e81000",
		16#2dbd# => X"e0ed3800",
		16#2dbe# => X"e4423800",
		16#2dbf# => X"13ffff96",
		16#2dc0# => X"e4223800",
		16#2dc1# => X"03fffff5",
		16#2dc2# => X"15000000",
		16#2dc3# => X"d4013808",
		16#2dc4# => X"a44300ff",
		16#2dc5# => X"bc220080",
		16#2dc6# => X"0c00002b",
		16#2dc7# => X"a4430100",
		16#2dc8# => X"9c400003",
		16#2dc9# => X"d4011810",
		16#2dca# => X"d401200c",
		16#2dcb# => X"d4011000",
		16#2dcc# => X"a8610000",
		16#2dcd# => X"07fffdf0",
		16#2dce# => X"15000000",
		16#2dcf# => X"9c210070",
		16#2dd0# => X"a84b0000",
		16#2dd1# => X"a86c0000",
		16#2dd2# => X"8521fffc",
		16#2dd3# => X"e1620004",
		16#2dd4# => X"e1830004",
		16#2dd5# => X"85c1ffe0",
		16#2dd6# => X"8441ffdc",
		16#2dd7# => X"8601ffe4",
		16#2dd8# => X"8641ffe8",
		16#2dd9# => X"8681ffec",
		16#2dda# => X"86c1fff0",
		16#2ddb# => X"8701fff4",
		16#2ddc# => X"44004800",
		16#2ddd# => X"8741fff8",
		16#2dde# => X"03ffff81",
		16#2ddf# => X"9d000000",
		16#2de0# => X"13ffff75",
		16#2de1# => X"9c400000",
		16#2de2# => X"03ffff75",
		16#2de3# => X"9c600000",
		16#2de4# => X"18600001",
		16#2de5# => X"bc050002",
		16#2de6# => X"13ffffe7",
		16#2de7# => X"a863877c",
		16#2de8# => X"8481002c",
		16#2de9# => X"84410018",
		16#2dea# => X"a86e0000",
		16#2deb# => X"e0441005",
		16#2dec# => X"e0801002",
		16#2ded# => X"e0441004",
		16#2dee# => X"b842005f",
		16#2def# => X"03ffffde",
		16#2df0# => X"d401102c",
		16#2df1# => X"bc220000",
		16#2df2# => X"13ffffd6",
		16#2df3# => X"e0a53004",
		16#2df4# => X"bc050000",
		16#2df5# => X"13ffffd3",
		16#2df6# => X"9ca30080",
		16#2df7# => X"e4851800",
		16#2df8# => X"10000003",
		16#2df9# => X"9cc00001",
		16#2dfa# => X"a8c20000",
		16#2dfb# => X"9ce0ff00",
		16#2dfc# => X"e0862000",
		16#2dfd# => X"03ffffcb",
		16#2dfe# => X"e0653803",
		16#2dff# => X"18600001",
		16#2e00# => X"bc020002",
		16#2e01# => X"13ffffcc",
		16#2e02# => X"a863877c",
		16#2e03# => X"84410018",
		16#2e04# => X"8481002c",
		16#2e05# => X"a8700000",
		16#2e06# => X"e0441005",
		16#2e07# => X"e0801002",
		16#2e08# => X"e0441004",
		16#2e09# => X"b842005f",
		16#2e0a# => X"03ffffc3",
		16#2e0b# => X"d4011018",
		16#2e0c# => X"d7e14ffc",
		16#2e0d# => X"d7e117f0",
		16#2e0e# => X"d7e177f4",
		16#2e0f# => X"d7e187f8",
		16#2e10# => X"9c21ffb8",
		16#2e11# => X"9dc10014",
		16#2e12# => X"d4011830",
		16#2e13# => X"d4012034",
		16#2e14# => X"9c610030",
		16#2e15# => X"d4012828",
		16#2e16# => X"d401302c",
		16#2e17# => X"07fffe5f",
		16#2e18# => X"a88e0000",
		16#2e19# => X"9c610028",
		16#2e1a# => X"07fffe5c",
		16#2e1b# => X"a8810000",
		16#2e1c# => X"84410014",
		16#2e1d# => X"bca20001",
		16#2e1e# => X"10000059",
		16#2e1f# => X"a86e0000",
		16#2e20# => X"84a10000",
		16#2e21# => X"bca50001",
		16#2e22# => X"10000055",
		16#2e23# => X"a8610000",
		16#2e24# => X"84810018",
		16#2e25# => X"84610004",
		16#2e26# => X"bc020004",
		16#2e27# => X"e0641805",
		16#2e28# => X"10000063",
		16#2e29# => X"d4011818",
		16#2e2a# => X"bc220002",
		16#2e2b# => X"0c000060",
		16#2e2c# => X"bc250004",
		16#2e2d# => X"0c000080",
		16#2e2e# => X"bc250002",
		16#2e2f# => X"0c00007a",
		16#2e30# => X"84410008",
		16#2e31# => X"8461001c",
		16#2e32# => X"84c10020",
		16#2e33# => X"e0431002",
		16#2e34# => X"8621000c",
		16#2e35# => X"d401101c",
		16#2e36# => X"84a10024",
		16#2e37# => X"e4513000",
		16#2e38# => X"0c00004b",
		16#2e39# => X"86e10010",
		16#2e3a# => X"e0652800",
		16#2e3b# => X"e4832800",
		16#2e3c# => X"0c000055",
		16#2e3d# => X"9c800001",
		16#2e3e# => X"e0c63000",
		16#2e3f# => X"9c42ffff",
		16#2e40# => X"e0c43000",
		16#2e41# => X"a8a30000",
		16#2e42# => X"d401101c",
		16#2e43# => X"9da0003d",
		16#2e44# => X"18401000",
		16#2e45# => X"9c600000",
		16#2e46# => X"9d600000",
		16#2e47# => X"9d800000",
		16#2e48# => X"baa2001f",
		16#2e49# => X"b9e30041",
		16#2e4a# => X"ba620041",
		16#2e4b# => X"9dadffff",
		16#2e4c# => X"e1f57804",
		16#2e4d# => X"a8f30000",
		16#2e4e# => X"e4513000",
		16#2e4f# => X"10000015",
		16#2e50# => X"a90f0000",
		16#2e51# => X"e1eb1004",
		16#2e52# => X"e2ac1804",
		16#2e53# => X"a84f0000",
		16#2e54# => X"e2668802",
		16#2e55# => X"e1e5b802",
		16#2e56# => X"e4313000",
		16#2e57# => X"10000005",
		16#2e58# => X"a8750000",
		16#2e59# => X"e4572800",
		16#2e5a# => X"1000000a",
		16#2e5b# => X"15000000",
		16#2e5c# => X"e44f2800",
		16#2e5d# => X"9cc00001",
		16#2e5e# => X"e1620004",
		16#2e5f# => X"e1830004",
		16#2e60# => X"10000003",
		16#2e61# => X"a8af0000",
		16#2e62# => X"9cc00000",
		16#2e63# => X"e0d33002",
		16#2e64# => X"e1e52800",
		16#2e65# => X"e0c63000",
		16#2e66# => X"e48f2800",
		16#2e67# => X"e0470004",
		16#2e68# => X"e0680004",
		16#2e69# => X"10000003",
		16#2e6a# => X"9e600001",
		16#2e6b# => X"9e600000",
		16#2e6c# => X"a8af0000",
		16#2e6d# => X"bc2d0000",
		16#2e6e# => X"13ffffda",
		16#2e6f# => X"e0d33000",
		16#2e70# => X"a46c00ff",
		16#2e71# => X"bc230080",
		16#2e72# => X"0c000026",
		16#2e73# => X"a88b0000",
		16#2e74# => X"a86e0000",
		16#2e75# => X"d4015820",
		16#2e76# => X"d4016024",
		16#2e77# => X"07fffd46",
		16#2e78# => X"15000000",
		16#2e79# => X"9c210048",
		16#2e7a# => X"a84b0000",
		16#2e7b# => X"a86c0000",
		16#2e7c# => X"8521fffc",
		16#2e7d# => X"e1620004",
		16#2e7e# => X"e1830004",
		16#2e7f# => X"85c1fff4",
		16#2e80# => X"8441fff0",
		16#2e81# => X"44004800",
		16#2e82# => X"8601fff8",
		16#2e83# => X"e4313000",
		16#2e84# => X"13ffffc0",
		16#2e85# => X"9da0003d",
		16#2e86# => X"e4572800",
		16#2e87# => X"0fffffbd",
		16#2e88# => X"e0652800",
		16#2e89# => X"03ffffb3",
		16#2e8a# => X"e4832800",
		16#2e8b# => X"18600001",
		16#2e8c# => X"e4022800",
		16#2e8d# => X"13ffffea",
		16#2e8e# => X"a863877c",
		16#2e8f# => X"03ffffe8",
		16#2e90# => X"a86e0000",
		16#2e91# => X"9c800000",
		16#2e92# => X"e0c63000",
		16#2e93# => X"9c42ffff",
		16#2e94# => X"e0c43000",
		16#2e95# => X"a8a30000",
		16#2e96# => X"03ffffad",
		16#2e97# => X"d401101c",
		16#2e98# => X"a46c0100",
		16#2e99# => X"bc230000",
		16#2e9a# => X"13ffffdb",
		16#2e9b# => X"a86e0000",
		16#2e9c# => X"e0c67804",
		16#2e9d# => X"bc060000",
		16#2e9e# => X"13ffffd7",
		16#2e9f# => X"15000000",
		16#2ea0# => X"9c6c0080",
		16#2ea1# => X"e4836000",
		16#2ea2# => X"10000003",
		16#2ea3# => X"9ca00001",
		16#2ea4# => X"a8ad0000",
		16#2ea5# => X"9c40ff00",
		16#2ea6# => X"e1652000",
		16#2ea7# => X"03ffffcd",
		16#2ea8# => X"e1831003",
		16#2ea9# => X"9c400004",
		16#2eaa# => X"a86e0000",
		16#2eab# => X"03ffffcc",
		16#2eac# => X"d4011014",
		16#2ead# => X"9c600000",
		16#2eae# => X"9c400000",
		16#2eaf# => X"d4011020",
		16#2eb0# => X"d4011824",
		16#2eb1# => X"9c600000",
		16#2eb2# => X"d401181c",
		16#2eb3# => X"03ffffc4",
		16#2eb4# => X"a86e0000",
		16#2eb5# => X"84a30000",
		16#2eb6# => X"9d600001",
		16#2eb7# => X"e4a55800",
		16#2eb8# => X"10000016",
		16#2eb9# => X"15000000",
		16#2eba# => X"84c40000",
		16#2ebb# => X"e4a65800",
		16#2ebc# => X"10000012",
		16#2ebd# => X"bc250004",
		16#2ebe# => X"0c000044",
		16#2ebf# => X"bc260004",
		16#2ec0# => X"0c000019",
		16#2ec1# => X"bc250002",
		16#2ec2# => X"0c000014",
		16#2ec3# => X"bc260002",
		16#2ec4# => X"0c00000c",
		16#2ec5# => X"15000000",
		16#2ec6# => X"84a30004",
		16#2ec7# => X"84c40004",
		16#2ec8# => X"e4053000",
		16#2ec9# => X"10000016",
		16#2eca# => X"15000000",
		16#2ecb# => X"bc050000",
		16#2ecc# => X"0c000008",
		16#2ecd# => X"15000000",
		16#2ece# => X"44004800",
		16#2ecf# => X"15000000",
		16#2ed0# => X"84630004",
		16#2ed1# => X"bc030000",
		16#2ed2# => X"13fffffc",
		16#2ed3# => X"15000000",
		16#2ed4# => X"44004800",
		16#2ed5# => X"9d60ffff",
		16#2ed6# => X"bc060002",
		16#2ed7# => X"13fffff7",
		16#2ed8# => X"9d600000",
		16#2ed9# => X"84640004",
		16#2eda# => X"bc030000",
		16#2edb# => X"13fffff3",
		16#2edc# => X"9d60ffff",
		16#2edd# => X"44004800",
		16#2ede# => X"9d600001",
		16#2edf# => X"84e30008",
		16#2ee0# => X"84c40008",
		16#2ee1# => X"e5a73000",
		16#2ee2# => X"0fffffea",
		16#2ee3# => X"bc050000",
		16#2ee4# => X"e5673000",
		16#2ee5# => X"0c000015",
		16#2ee6# => X"bc050000",
		16#2ee7# => X"84c3000c",
		16#2ee8# => X"84e4000c",
		16#2ee9# => X"84630010",
		16#2eea# => X"e4463800",
		16#2eeb# => X"10000013",
		16#2eec# => X"84840010",
		16#2eed# => X"e4263800",
		16#2eee# => X"10000005",
		16#2eef# => X"e4473000",
		16#2ef0# => X"e4432000",
		16#2ef1# => X"1000000d",
		16#2ef2# => X"e4473000",
		16#2ef3# => X"10000007",
		16#2ef4# => X"bc050000",
		16#2ef5# => X"e4273000",
		16#2ef6# => X"1000000a",
		16#2ef7# => X"e4441800",
		16#2ef8# => X"0c000008",
		16#2ef9# => X"bc050000",
		16#2efa# => X"0fffffe3",
		16#2efb# => X"9d60ffff",
		16#2efc# => X"44004800",
		16#2efd# => X"15000000",
		16#2efe# => X"03ffffcd",
		16#2eff# => X"9d600001",
		16#2f00# => X"44004800",
		16#2f01# => X"9d600000",
		16#2f02# => X"13ffffce",
		16#2f03# => X"15000000",
		16#2f04# => X"85640004",
		16#2f05# => X"84630004",
		16#2f06# => X"44004800",
		16#2f07# => X"e16b1802",
		16#2f08# => X"d7e14ffc",
		16#2f09# => X"d7e117f4",
		16#2f0a# => X"d7e177f8",
		16#2f0b# => X"9c21ffbc",
		16#2f0c# => X"9dc10014",
		16#2f0d# => X"d4011830",
		16#2f0e# => X"d4012034",
		16#2f0f# => X"9c610030",
		16#2f10# => X"d4012828",
		16#2f11# => X"d401302c",
		16#2f12# => X"07fffd64",
		16#2f13# => X"a88e0000",
		16#2f14# => X"9c610028",
		16#2f15# => X"07fffd61",
		16#2f16# => X"a8810000",
		16#2f17# => X"a86e0000",
		16#2f18# => X"07ffff9d",
		16#2f19# => X"a8810000",
		16#2f1a# => X"9c210044",
		16#2f1b# => X"8521fffc",
		16#2f1c# => X"8441fff4",
		16#2f1d# => X"44004800",
		16#2f1e# => X"85c1fff8",
		16#2f1f# => X"d7e14ffc",
		16#2f20# => X"d7e177f8",
		16#2f21# => X"d7e117f4",
		16#2f22# => X"9c21ffbc",
		16#2f23# => X"9dc10014",
		16#2f24# => X"d4011830",
		16#2f25# => X"d4012034",
		16#2f26# => X"9c610030",
		16#2f27# => X"d4012828",
		16#2f28# => X"d401302c",
		16#2f29# => X"07fffd4d",
		16#2f2a# => X"a88e0000",
		16#2f2b# => X"9c610028",
		16#2f2c# => X"07fffd4a",
		16#2f2d# => X"a8810000",
		16#2f2e# => X"9d600001",
		16#2f2f# => X"84610014",
		16#2f30# => X"e4a35800",
		16#2f31# => X"10000007",
		16#2f32# => X"84610000",
		16#2f33# => X"e4a35800",
		16#2f34# => X"10000004",
		16#2f35# => X"a86e0000",
		16#2f36# => X"07ffff7f",
		16#2f37# => X"a8810000",
		16#2f38# => X"9c210044",
		16#2f39# => X"8521fffc",
		16#2f3a# => X"8441fff4",
		16#2f3b# => X"44004800",
		16#2f3c# => X"85c1fff8",
		16#2f3d# => X"d7e14ffc",
		16#2f3e# => X"d7e177f8",
		16#2f3f# => X"d7e117f4",
		16#2f40# => X"9c21ffbc",
		16#2f41# => X"9dc10014",
		16#2f42# => X"d4011830",
		16#2f43# => X"d4012034",
		16#2f44# => X"9c610030",
		16#2f45# => X"d4012828",
		16#2f46# => X"d401302c",
		16#2f47# => X"07fffd2f",
		16#2f48# => X"a88e0000",
		16#2f49# => X"9c610028",
		16#2f4a# => X"07fffd2c",
		16#2f4b# => X"a8810000",
		16#2f4c# => X"9d600001",
		16#2f4d# => X"84610014",
		16#2f4e# => X"e4a35800",
		16#2f4f# => X"10000007",
		16#2f50# => X"84610000",
		16#2f51# => X"e4a35800",
		16#2f52# => X"10000004",
		16#2f53# => X"a86e0000",
		16#2f54# => X"07ffff61",
		16#2f55# => X"a8810000",
		16#2f56# => X"9c210044",
		16#2f57# => X"8521fffc",
		16#2f58# => X"8441fff4",
		16#2f59# => X"44004800",
		16#2f5a# => X"85c1fff8",
		16#2f5b# => X"d7e14ffc",
		16#2f5c# => X"d7e177f8",
		16#2f5d# => X"d7e117f4",
		16#2f5e# => X"9c21ffbc",
		16#2f5f# => X"9dc10014",
		16#2f60# => X"d4011830",
		16#2f61# => X"d4012034",
		16#2f62# => X"9c610030",
		16#2f63# => X"d4012828",
		16#2f64# => X"d401302c",
		16#2f65# => X"07fffd11",
		16#2f66# => X"a88e0000",
		16#2f67# => X"9c610028",
		16#2f68# => X"07fffd0e",
		16#2f69# => X"a8810000",
		16#2f6a# => X"84610014",
		16#2f6b# => X"bca30001",
		16#2f6c# => X"10000008",
		16#2f6d# => X"9d60ffff",
		16#2f6e# => X"84610000",
		16#2f6f# => X"bca30001",
		16#2f70# => X"10000004",
		16#2f71# => X"a86e0000",
		16#2f72# => X"07ffff43",
		16#2f73# => X"a8810000",
		16#2f74# => X"9c210044",
		16#2f75# => X"8521fffc",
		16#2f76# => X"8441fff4",
		16#2f77# => X"44004800",
		16#2f78# => X"85c1fff8",
		16#2f79# => X"d7e14ffc",
		16#2f7a# => X"d7e177f8",
		16#2f7b# => X"d7e117f4",
		16#2f7c# => X"9c21ffbc",
		16#2f7d# => X"9dc10014",
		16#2f7e# => X"d4011830",
		16#2f7f# => X"d4012034",
		16#2f80# => X"9c610030",
		16#2f81# => X"d4012828",
		16#2f82# => X"d401302c",
		16#2f83# => X"07fffcf3",
		16#2f84# => X"a88e0000",
		16#2f85# => X"9c610028",
		16#2f86# => X"07fffcf0",
		16#2f87# => X"a8810000",
		16#2f88# => X"84610014",
		16#2f89# => X"bca30001",
		16#2f8a# => X"10000008",
		16#2f8b# => X"9d60ffff",
		16#2f8c# => X"84610000",
		16#2f8d# => X"bca30001",
		16#2f8e# => X"10000004",
		16#2f8f# => X"a86e0000",
		16#2f90# => X"07ffff25",
		16#2f91# => X"a8810000",
		16#2f92# => X"9c210044",
		16#2f93# => X"8521fffc",
		16#2f94# => X"8441fff4",
		16#2f95# => X"44004800",
		16#2f96# => X"85c1fff8",
		16#2f97# => X"d7e14ffc",
		16#2f98# => X"d7e177f8",
		16#2f99# => X"d7e117f4",
		16#2f9a# => X"9c21ffbc",
		16#2f9b# => X"9dc10014",
		16#2f9c# => X"d4011830",
		16#2f9d# => X"d4012034",
		16#2f9e# => X"9c610030",
		16#2f9f# => X"d4012828",
		16#2fa0# => X"d401302c",
		16#2fa1# => X"07fffcd5",
		16#2fa2# => X"a88e0000",
		16#2fa3# => X"9c610028",
		16#2fa4# => X"07fffcd2",
		16#2fa5# => X"a8810000",
		16#2fa6# => X"9d600001",
		16#2fa7# => X"84610014",
		16#2fa8# => X"e4a35800",
		16#2fa9# => X"10000007",
		16#2faa# => X"84610000",
		16#2fab# => X"e4a35800",
		16#2fac# => X"10000004",
		16#2fad# => X"a86e0000",
		16#2fae# => X"07ffff07",
		16#2faf# => X"a8810000",
		16#2fb0# => X"9c210044",
		16#2fb1# => X"8521fffc",
		16#2fb2# => X"8441fff4",
		16#2fb3# => X"44004800",
		16#2fb4# => X"85c1fff8",
		16#2fb5# => X"d7e14ffc",
		16#2fb6# => X"d7e177f8",
		16#2fb7# => X"d7e117f4",
		16#2fb8# => X"9c21ffbc",
		16#2fb9# => X"9dc10014",
		16#2fba# => X"d4011830",
		16#2fbb# => X"d4012034",
		16#2fbc# => X"9c610030",
		16#2fbd# => X"d4012828",
		16#2fbe# => X"d401302c",
		16#2fbf# => X"07fffcb7",
		16#2fc0# => X"a88e0000",
		16#2fc1# => X"9c610028",
		16#2fc2# => X"07fffcb4",
		16#2fc3# => X"a8810000",
		16#2fc4# => X"9d600001",
		16#2fc5# => X"84610014",
		16#2fc6# => X"e4a35800",
		16#2fc7# => X"10000007",
		16#2fc8# => X"84610000",
		16#2fc9# => X"e4a35800",
		16#2fca# => X"10000004",
		16#2fcb# => X"a86e0000",
		16#2fcc# => X"07fffee9",
		16#2fcd# => X"a8810000",
		16#2fce# => X"9c210044",
		16#2fcf# => X"8521fffc",
		16#2fd0# => X"8441fff4",
		16#2fd1# => X"44004800",
		16#2fd2# => X"85c1fff8",
		16#2fd3# => X"d7e14ffc",
		16#2fd4# => X"9c21ffc4",
		16#2fd5# => X"d4011830",
		16#2fd6# => X"d4012034",
		16#2fd7# => X"9c610030",
		16#2fd8# => X"d4012828",
		16#2fd9# => X"d401302c",
		16#2fda# => X"07fffc9c",
		16#2fdb# => X"9c810014",
		16#2fdc# => X"9c610028",
		16#2fdd# => X"07fffc99",
		16#2fde# => X"a8810000",
		16#2fdf# => X"9d600001",
		16#2fe0# => X"84610014",
		16#2fe1# => X"e4a35800",
		16#2fe2# => X"10000005",
		16#2fe3# => X"84610000",
		16#2fe4# => X"e4a35800",
		16#2fe5# => X"0c000006",
		16#2fe6# => X"15000000",
		16#2fe7# => X"9c21003c",
		16#2fe8# => X"8521fffc",
		16#2fe9# => X"44004800",
		16#2fea# => X"15000000",
		16#2feb# => X"9c21003c",
		16#2fec# => X"8521fffc",
		16#2fed# => X"44004800",
		16#2fee# => X"9d600000",
		16#2fef# => X"b883005f",
		16#2ff0# => X"d7e117f8",
		16#2ff1# => X"d7e14ffc",
		16#2ff2# => X"9c400003",
		16#2ff3# => X"9c21ffe4",
		16#2ff4# => X"bc230000",
		16#2ff5# => X"d4011000",
		16#2ff6# => X"1000000a",
		16#2ff7# => X"d4012004",
		16#2ff8# => X"9c400002",
		16#2ff9# => X"d4011000",
		16#2ffa# => X"07fffbc3",
		16#2ffb# => X"a8610000",
		16#2ffc# => X"9c21001c",
		16#2ffd# => X"8521fffc",
		16#2ffe# => X"44004800",
		16#2fff# => X"8441fff8",
		16#3000# => X"a8430000",
		16#3001# => X"9c60003c",
		16#3002# => X"bc040000",
		16#3003# => X"0c000015",
		16#3004# => X"d4011808",
		16#3005# => X"9c800000",
		16#3006# => X"a8620000",
		16#3007# => X"d401200c",
		16#3008# => X"04000134",
		16#3009# => X"d4011010",
		16#300a# => X"9c8b001d",
		16#300b# => X"bda40000",
		16#300c# => X"13ffffee",
		16#300d# => X"9d6bfffd",
		16#300e# => X"bd8b0000",
		16#300f# => X"1000000f",
		16#3010# => X"e1625808",
		16#3011# => X"9c400000",
		16#3012# => X"d401580c",
		16#3013# => X"d4011010",
		16#3014# => X"9c40003c",
		16#3015# => X"e0822002",
		16#3016# => X"03ffffe4",
		16#3017# => X"d4012008",
		16#3018# => X"18608000",
		16#3019# => X"e4021800",
		16#301a# => X"1000000c",
		16#301b# => X"1960c1e0",
		16#301c# => X"03ffffe9",
		16#301d# => X"e0401002",
		16#301e# => X"9ca0001f",
		16#301f# => X"b8620041",
		16#3020# => X"e0a52002",
		16#3021# => X"e0422008",
		16#3022# => X"e0a32848",
		16#3023# => X"d4011010",
		16#3024# => X"03fffff0",
		16#3025# => X"d401280c",
		16#3026# => X"03ffffd6",
		16#3027# => X"9d800000",
		16#3028# => X"d7e117f8",
		16#3029# => X"9c800000",
		16#302a# => X"d7e14ffc",
		16#302b# => X"9c21ffe4",
		16#302c# => X"a8430000",
		16#302d# => X"e4232000",
		16#302e# => X"0c000023",
		16#302f# => X"d4012004",
		16#3030# => X"9c800003",
		16#3031# => X"9ca00000",
		16#3032# => X"d4012000",
		16#3033# => X"9c80003c",
		16#3034# => X"d4011810",
		16#3035# => X"d4012008",
		16#3036# => X"04000106",
		16#3037# => X"d401280c",
		16#3038# => X"9c6b001d",
		16#3039# => X"bd630000",
		16#303a# => X"0c00001a",
		16#303b# => X"bc030000",
		16#303c# => X"1000000b",
		16#303d# => X"9d6bfffd",
		16#303e# => X"bd8b0000",
		16#303f# => X"1000002a",
		16#3040# => X"e1625808",
		16#3041# => X"9c400000",
		16#3042# => X"d401580c",
		16#3043# => X"d4011010",
		16#3044# => X"9c40003c",
		16#3045# => X"e0621802",
		16#3046# => X"d4011808",
		16#3047# => X"07fffb76",
		16#3048# => X"a8610000",
		16#3049# => X"9c21001c",
		16#304a# => X"a84b0000",
		16#304b# => X"a86c0000",
		16#304c# => X"8521fffc",
		16#304d# => X"e1620004",
		16#304e# => X"e1830004",
		16#304f# => X"44004800",
		16#3050# => X"8441fff8",
		16#3051# => X"9c400002",
		16#3052# => X"03fffff5",
		16#3053# => X"d4011000",
		16#3054# => X"e0801802",
		16#3055# => X"9cc4ffe0",
		16#3056# => X"bd860000",
		16#3057# => X"1000001a",
		16#3058# => X"9ca00000",
		16#3059# => X"9ca5ffff",
		16#305a# => X"e0822048",
		16#305b# => X"e0a51003",
		16#305c# => X"b8c6009f",
		16#305d# => X"e0402802",
		16#305e# => X"e0a22804",
		16#305f# => X"e0843003",
		16#3060# => X"b845005f",
		16#3061# => X"9ca0003c",
		16#3062# => X"e0422004",
		16#3063# => X"e0651802",
		16#3064# => X"9ca00000",
		16#3065# => X"d4011808",
		16#3066# => X"d401280c",
		16#3067# => X"03ffffe0",
		16#3068# => X"d4011010",
		16#3069# => X"9c80001f",
		16#306a# => X"b8a20041",
		16#306b# => X"e0841802",
		16#306c# => X"e0421808",
		16#306d# => X"e0852048",
		16#306e# => X"d4011010",
		16#306f# => X"03ffffd5",
		16#3070# => X"d401200c",
		16#3071# => X"9ca00001",
		16#3072# => X"03ffffe7",
		16#3073# => X"e0a52008",
		16#3074# => X"d7e14ffc",
		16#3075# => X"9c21ffe0",
		16#3076# => X"d4011814",
		16#3077# => X"d4012018",
		16#3078# => X"9c610014",
		16#3079# => X"07fffbfd",
		16#307a# => X"a8810000",
		16#307b# => X"84610000",
		16#307c# => X"bc030002",
		16#307d# => X"10000018",
		16#307e# => X"9d600000",
		16#307f# => X"bca30001",
		16#3080# => X"10000015",
		16#3081# => X"bc230004",
		16#3082# => X"0c000020",
		16#3083# => X"84610008",
		16#3084# => X"bd830000",
		16#3085# => X"10000010",
		16#3086# => X"bda3001e",
		16#3087# => X"0c000012",
		16#3088# => X"9d60003c",
		16#3089# => X"e06b1802",
		16#308a# => X"9c83ffe0",
		16#308b# => X"bd840000",
		16#308c# => X"1000001e",
		16#308d# => X"84a1000c",
		16#308e# => X"8561000c",
		16#308f# => X"e16b2048",
		16#3090# => X"84610004",
		16#3091# => X"bc030000",
		16#3092# => X"10000003",
		16#3093# => X"15000000",
		16#3094# => X"e1605802",
		16#3095# => X"9c210020",
		16#3096# => X"8521fffc",
		16#3097# => X"44004800",
		16#3098# => X"15000000",
		16#3099# => X"84610004",
		16#309a# => X"bc030000",
		16#309b# => X"0c00000b",
		16#309c# => X"15000000",
		16#309d# => X"9c210020",
		16#309e# => X"19607fff",
		16#309f# => X"8521fffc",
		16#30a0# => X"44004800",
		16#30a1# => X"a96bffff",
		16#30a2# => X"84610004",
		16#30a3# => X"e4035800",
		16#30a4# => X"13fffff9",
		16#30a5# => X"15000000",
		16#30a6# => X"9c210020",
		16#30a7# => X"8521fffc",
		16#30a8# => X"44004800",
		16#30a9# => X"19608000",
		16#30aa# => X"9c80001f",
		16#30ab# => X"b8a50001",
		16#30ac# => X"e0841802",
		16#30ad# => X"85610010",
		16#30ae# => X"e0852008",
		16#30af# => X"e16b1848",
		16#30b0# => X"03ffffe0",
		16#30b1# => X"e1645804",
		16#30b2# => X"d7e14ffc",
		16#30b3# => X"d7e117f8",
		16#30b4# => X"9c21ffdc",
		16#30b5# => X"d4011814",
		16#30b6# => X"d4012018",
		16#30b7# => X"9c610014",
		16#30b8# => X"07fffbbe",
		16#30b9# => X"a8810000",
		16#30ba# => X"84810004",
		16#30bb# => X"a8610000",
		16#30bc# => X"e0402002",
		16#30bd# => X"e0422004",
		16#30be# => X"ac42ffff",
		16#30bf# => X"b842005f",
		16#30c0# => X"07fffafd",
		16#30c1# => X"d4011004",
		16#30c2# => X"9c210024",
		16#30c3# => X"a84b0000",
		16#30c4# => X"a86c0000",
		16#30c5# => X"8521fffc",
		16#30c6# => X"e1620004",
		16#30c7# => X"e1830004",
		16#30c8# => X"44004800",
		16#30c9# => X"8441fff8",
		16#30ca# => X"d7e14ffc",
		16#30cb# => X"d7e117f8",
		16#30cc# => X"9c21ffe4",
		16#30cd# => X"d4011800",
		16#30ce# => X"d4012004",
		16#30cf# => X"d4012808",
		16#30d0# => X"d401300c",
		16#30d1# => X"d4013810",
		16#30d2# => X"07fffaeb",
		16#30d3# => X"a8610000",
		16#30d4# => X"9c21001c",
		16#30d5# => X"a84b0000",
		16#30d6# => X"a86c0000",
		16#30d7# => X"8521fffc",
		16#30d8# => X"e1620004",
		16#30d9# => X"e1830004",
		16#30da# => X"44004800",
		16#30db# => X"8441fff8",
		16#30dc# => X"d7e117f8",
		16#30dd# => X"d7e14ffc",
		16#30de# => X"9c21ffdc",
		16#30df# => X"18403fff",
		16#30e0# => X"d4011814",
		16#30e1# => X"d4012018",
		16#30e2# => X"9c610014",
		16#30e3# => X"a8810000",
		16#30e4# => X"07fffb92",
		16#30e5# => X"a842ffff",
		16#30e6# => X"84610010",
		16#30e7# => X"84c1000c",
		16#30e8# => X"b883005e",
		16#30e9# => X"b8c60002",
		16#30ea# => X"e0631003",
		16#30eb# => X"bc030000",
		16#30ec# => X"10000003",
		16#30ed# => X"e0c62004",
		16#30ee# => X"a8c60001",
		16#30ef# => X"84610000",
		16#30f0# => X"84810004",
		16#30f1# => X"07fff98b",
		16#30f2# => X"84a10008",
		16#30f3# => X"9c210024",
		16#30f4# => X"8521fffc",
		16#30f5# => X"44004800",
		16#30f6# => X"8441fff8",
		16#30f7# => X"a4e4ffff",
		16#30f8# => X"b9040050",
		16#30f9# => X"a566ffff",
		16#30fa# => X"b9860050",
		16#30fb# => X"e1ab3b06",
		16#30fc# => X"e16b4306",
		16#30fd# => X"e0ec3b06",
		16#30fe# => X"b9ed0050",
		16#30ff# => X"e0eb3800",
		16#3100# => X"d7e117fc",
		16#3101# => X"e0e77800",
		16#3102# => X"9c21fffc",
		16#3103# => X"e4ab3800",
		16#3104# => X"10000004",
		16#3105# => X"e10c4306",
		16#3106# => X"18400001",
		16#3107# => X"e1081000",
		16#3108# => X"e0c61b06",
		16#3109# => X"e0842b06",
		16#310a# => X"b8670050",
		16#310b# => X"b8e70010",
		16#310c# => X"a5adffff",
		16#310d# => X"e1081800",
		16#310e# => X"e1643000",
		16#310f# => X"9c210004",
		16#3110# => X"e1876800",
		16#3111# => X"e16b4000",
		16#3112# => X"44004800",
		16#3113# => X"8441fffc",
		16#3114# => X"bc050000",
		16#3115# => X"1000000b",
		16#3116# => X"9cc00020",
		16#3117# => X"e0c62802",
		16#3118# => X"bd460000",
		16#3119# => X"0c00000a",
		16#311a# => X"15000000",
		16#311b# => X"e0c33008",
		16#311c# => X"e0842848",
		16#311d# => X"e0a32848",
		16#311e# => X"e0862004",
		16#311f# => X"a8650000",
		16#3120# => X"a9630000",
		16#3121# => X"44004800",
		16#3122# => X"a9840000",
		16#3123# => X"e0803002",
		16#3124# => X"9ca00000",
		16#3125# => X"e0832048",
		16#3126# => X"03fffffa",
		16#3127# => X"a8650000",
		16#3128# => X"bc050000",
		16#3129# => X"1000000b",
		16#312a# => X"9cc00020",
		16#312b# => X"e0c62802",
		16#312c# => X"bd460000",
		16#312d# => X"0c00000a",
		16#312e# => X"15000000",
		16#312f# => X"e0c43048",
		16#3130# => X"e0632808",
		16#3131# => X"e0a42808",
		16#3132# => X"e0661804",
		16#3133# => X"a8850000",
		16#3134# => X"a9630000",
		16#3135# => X"44004800",
		16#3136# => X"a9840000",
		16#3137# => X"e0603002",
		16#3138# => X"9ca00000",
		16#3139# => X"e0641808",
		16#313a# => X"03fffffa",
		16#313b# => X"a8850000",
		16#313c# => X"d7e117fc",
		16#313d# => X"a840ffff",
		16#313e# => X"e4431000",
		16#313f# => X"10000010",
		16#3140# => X"9c21fffc",
		16#3141# => X"bc4300ff",
		16#3142# => X"0c000018",
		16#3143# => X"9c800020",
		16#3144# => X"9c800018",
		16#3145# => X"9ca00008",
		16#3146# => X"18400001",
		16#3147# => X"e0632848",
		16#3148# => X"a8428790",
		16#3149# => X"9c210004",
		16#314a# => X"e0631000",
		16#314b# => X"8441fffc",
		16#314c# => X"8d630000",
		16#314d# => X"44004800",
		16#314e# => X"e1645802",
		16#314f# => X"184000ff",
		16#3150# => X"a842ffff",
		16#3151# => X"e4431000",
		16#3152# => X"10000005",
		16#3153# => X"15000000",
		16#3154# => X"9c800010",
		16#3155# => X"03fffff1",
		16#3156# => X"a8a40000",
		16#3157# => X"9c800008",
		16#3158# => X"03ffffee",
		16#3159# => X"9ca00018",
		16#315a# => X"03ffffec",
		16#315b# => X"9ca00000",
		16#315c# => X"d7e14ffc",
		16#315d# => X"9c21fffc",
		16#315e# => X"a8830000",
		16#315f# => X"9c210004",
		16#3160# => X"9c600000",
		16#3161# => X"8521fffc",
		16#3162# => X"a8a30000",
		16#3163# => X"00000e88",
		16#3164# => X"a8c30000",
		16#3165# => X"d7e117f8",
		16#3166# => X"d7e14ffc",
		16#3167# => X"9c800000",
		16#3168# => X"9c21fff8",
		16#3169# => X"04000ed3",
		16#316a# => X"a8430000",
		16#316b# => X"18800001",
		16#316c# => X"a8848890",
		16#316d# => X"84840000",
		16#316e# => X"84a4003c",
		16#316f# => X"bc050000",
		16#3170# => X"10000004",
		16#3171# => X"15000000",
		16#3172# => X"48002800",
		16#3173# => X"a8640000",
		16#3174# => X"04002c48",
		16#3175# => X"a8620000",
		16#3176# => X"a8830000",
		16#3177# => X"18600001",
		16#3178# => X"d7e14ffc",
		16#3179# => X"a863ade4",
		16#317a# => X"9c21fffc",
		16#317b# => X"84630000",
		16#317c# => X"9c210004",
		16#317d# => X"8521fffc",
		16#317e# => X"0000000c",
		16#317f# => X"15000000",
		16#3180# => X"a8830000",
		16#3181# => X"18600001",
		16#3182# => X"d7e14ffc",
		16#3183# => X"a863ade4",
		16#3184# => X"9c21fffc",
		16#3185# => X"84630000",
		16#3186# => X"9c210004",
		16#3187# => X"8521fffc",
		16#3188# => X"00001927",
		16#3189# => X"15000000",
		16#318a# => X"d7e177dc",
		16#318b# => X"d7e187e0",
		16#318c# => X"d7e14ffc",
		16#318d# => X"d7e117d8",
		16#318e# => X"d7e197e4",
		16#318f# => X"d7e1a7e8",
		16#3190# => X"d7e1b7ec",
		16#3191# => X"d7e1c7f0",
		16#3192# => X"d7e1d7f4",
		16#3193# => X"d7e1e7f8",
		16#3194# => X"9dc4000b",
		16#3195# => X"9c21ffd8",
		16#3196# => X"bcae0016",
		16#3197# => X"10000036",
		16#3198# => X"aa030000",
		16#3199# => X"9c40fff8",
		16#319a# => X"e1ce1003",
		16#319b# => X"b86e005f",
		16#319c# => X"e48e2000",
		16#319d# => X"10000003",
		16#319e# => X"9c400001",
		16#319f# => X"9c400000",
		16#31a0# => X"a44200ff",
		16#31a1# => X"bc220000",
		16#31a2# => X"100000b3",
		16#31a3# => X"bc030000",
		16#31a4# => X"0c0000b2",
		16#31a5# => X"9c40000c",
		16#31a6# => X"04000234",
		16#31a7# => X"a8700000",
		16#31a8# => X"bc4e01f7",
		16#31a9# => X"10000027",
		16#31aa# => X"b8ee0049",
		16#31ab# => X"18800001",
		16#31ac# => X"b8ee0043",
		16#31ad# => X"a884b20c",
		16#31ae# => X"e06e2000",
		16#31af# => X"8443000c",
		16#31b0# => X"e4221800",
		16#31b1# => X"0c00018e",
		16#31b2# => X"aa440000",
		16#31b3# => X"84820004",
		16#31b4# => X"9ca0fffc",
		16#31b5# => X"8462000c",
		16#31b6# => X"e0842803",
		16#31b7# => X"84c20008",
		16#31b8# => X"e0822000",
		16#31b9# => X"d406180c",
		16#31ba# => X"84a40004",
		16#31bb# => X"d4033008",
		16#31bc# => X"a8a50001",
		16#31bd# => X"a8700000",
		16#31be# => X"0400021e",
		16#31bf# => X"d4042804",
		16#31c0# => X"9d620008",
		16#31c1# => X"9c210028",
		16#31c2# => X"8521fffc",
		16#31c3# => X"8441ffd8",
		16#31c4# => X"85c1ffdc",
		16#31c5# => X"8601ffe0",
		16#31c6# => X"8641ffe4",
		16#31c7# => X"8681ffe8",
		16#31c8# => X"86c1ffec",
		16#31c9# => X"8701fff0",
		16#31ca# => X"8741fff4",
		16#31cb# => X"44004800",
		16#31cc# => X"8781fff8",
		16#31cd# => X"9c600000",
		16#31ce# => X"03ffffce",
		16#31cf# => X"9dc00010",
		16#31d0# => X"bc270000",
		16#31d1# => X"0c000088",
		16#31d2# => X"bc470004",
		16#31d3# => X"10000155",
		16#31d4# => X"bc470014",
		16#31d5# => X"b8ee0046",
		16#31d6# => X"9ce70038",
		16#31d7# => X"b8670003",
		16#31d8# => X"19600001",
		16#31d9# => X"a96bb20c",
		16#31da# => X"e0635800",
		16#31db# => X"8443000c",
		16#31dc# => X"e4031000",
		16#31dd# => X"10000019",
		16#31de# => X"aa4b0000",
		16#31df# => X"9ca0fffc",
		16#31e0# => X"84820004",
		16#31e1# => X"e0842803",
		16#31e2# => X"e0a47002",
		16#31e3# => X"bd45000f",
		16#31e4# => X"100000b9",
		16#31e5# => X"bd650000",
		16#31e6# => X"0c00000c",
		16#31e7# => X"15000000",
		16#31e8# => X"000000b8",
		16#31e9# => X"e0822000",
		16#31ea# => X"84820004",
		16#31eb# => X"e0845803",
		16#31ec# => X"e0a47002",
		16#31ed# => X"bda5000f",
		16#31ee# => X"0c0000af",
		16#31ef# => X"bd850000",
		16#31f0# => X"0c0000af",
		16#31f1# => X"15000000",
		16#31f2# => X"8442000c",
		16#31f3# => X"e4231000",
		16#31f4# => X"13fffff6",
		16#31f5# => X"9d60fffc",
		16#31f6# => X"9ce70001",
		16#31f7# => X"18c00001",
		16#31f8# => X"a8c6b214",
		16#31f9# => X"84460008",
		16#31fa# => X"e4261000",
		16#31fb# => X"0c00007f",
		16#31fc# => X"9c60fffc",
		16#31fd# => X"84820004",
		16#31fe# => X"e0841803",
		16#31ff# => X"e0647002",
		16#3200# => X"bda3000f",
		16#3201# => X"0c00012f",
		16#3202# => X"bd830000",
		16#3203# => X"d406300c",
		16#3204# => X"0c0000a7",
		16#3205# => X"d4063008",
		16#3206# => X"bc4401ff",
		16#3207# => X"10000055",
		16#3208# => X"b8640049",
		16#3209# => X"b8640043",
		16#320a# => X"9d000001",
		16#320b# => X"84920004",
		16#320c# => X"b8a30082",
		16#320d# => X"b8630003",
		16#320e# => X"e1082808",
		16#320f# => X"18a00001",
		16#3210# => X"a8a5b20c",
		16#3211# => X"e0882004",
		16#3212# => X"e0632800",
		16#3213# => X"d4122004",
		16#3214# => X"84a30008",
		16#3215# => X"d402180c",
		16#3216# => X"d4022808",
		16#3217# => X"d4031008",
		16#3218# => X"d405100c",
		16#3219# => X"b8470082",
		16#321a# => X"9c600001",
		16#321b# => X"e0631008",
		16#321c# => X"e4432000",
		16#321d# => X"10000064",
		16#321e# => X"e0441803",
		16#321f# => X"bc220000",
		16#3220# => X"1000000d",
		16#3221# => X"9c40fffc",
		16#3222# => X"e0631800",
		16#3223# => X"e0e71003",
		16#3224# => X"e0441803",
		16#3225# => X"bc220000",
		16#3226# => X"10000007",
		16#3227# => X"9ce70004",
		16#3228# => X"e0631800",
		16#3229# => X"e0432003",
		16#322a# => X"bc020000",
		16#322b# => X"13fffffd",
		16#322c# => X"9ce70004",
		16#322d# => X"18800001",
		16#322e# => X"b9870003",
		16#322f# => X"a884b20c",
		16#3230# => X"a9670000",
		16#3231# => X"e18c2000",
		16#3232# => X"a90c0000",
		16#3233# => X"8448000c",
		16#3234# => X"e4081000",
		16#3235# => X"10000019",
		16#3236# => X"9c80fffc",
		16#3237# => X"84a20004",
		16#3238# => X"e0a52003",
		16#3239# => X"e0857002",
		16#323a# => X"bd44000f",
		16#323b# => X"1000010b",
		16#323c# => X"bd640000",
		16#323d# => X"0c00000d",
		16#323e# => X"15000000",
		16#323f# => X"0000011b",
		16#3240# => X"e0a22800",
		16#3241# => X"9c80fffc",
		16#3242# => X"84a20004",
		16#3243# => X"e0a52003",
		16#3244# => X"e0857002",
		16#3245# => X"bda4000f",
		16#3246# => X"0c000100",
		16#3247# => X"bd840000",
		16#3248# => X"0c000111",
		16#3249# => X"15000000",
		16#324a# => X"8442000c",
		16#324b# => X"e4281000",
		16#324c# => X"13fffff5",
		16#324d# => X"15000000",
		16#324e# => X"9d6b0001",
		16#324f# => X"a44b0003",
		16#3250# => X"bc220000",
		16#3251# => X"0c000142",
		16#3252# => X"9d080008",
		16#3253# => X"03ffffe1",
		16#3254# => X"8448000c",
		16#3255# => X"9c40000c",
		16#3256# => X"9d600000",
		16#3257# => X"03ffff6a",
		16#3258# => X"d4101000",
		16#3259# => X"b8ee0043",
		16#325a# => X"03ffff7e",
		16#325b# => X"b8670003",
		16#325c# => X"bc430004",
		16#325d# => X"1000010b",
		16#325e# => X"bc430014",
		16#325f# => X"b9040046",
		16#3260# => X"9d080038",
		16#3261# => X"19600001",
		16#3262# => X"b8a80003",
		16#3263# => X"a96bb20c",
		16#3264# => X"e0a55800",
		16#3265# => X"84650008",
		16#3266# => X"e4032800",
		16#3267# => X"0c000008",
		16#3268# => X"b9080082",
		16#3269# => X"00000114",
		16#326a# => X"9c800001",
		16#326b# => X"84630008",
		16#326c# => X"e4051800",
		16#326d# => X"10000008",
		16#326e# => X"15000000",
		16#326f# => X"85030004",
		16#3270# => X"9d60fffc",
		16#3271# => X"e1085803",
		16#3272# => X"e4844000",
		16#3273# => X"13fffff8",
		16#3274# => X"15000000",
		16#3275# => X"8483000c",
		16#3276# => X"d402200c",
		16#3277# => X"d4021808",
		16#3278# => X"d4041008",
		16#3279# => X"d403100c",
		16#327a# => X"b8470082",
		16#327b# => X"9c600001",
		16#327c# => X"84920004",
		16#327d# => X"e0631008",
		16#327e# => X"e4432000",
		16#327f# => X"0fffffa0",
		16#3280# => X"e0441803",
		16#3281# => X"84520008",
		16#3282# => X"9ca0fffc",
		16#3283# => X"86820004",
		16#3284# => X"e2942803",
		16#3285# => X"e0747002",
		16#3286# => X"bda3000f",
		16#3287# => X"10000003",
		16#3288# => X"9c800001",
		16#3289# => X"9c800000",
		16#328a# => X"a48400ff",
		16#328b# => X"bc240000",
		16#328c# => X"10000027",
		16#328d# => X"e44ea000",
		16#328e# => X"0c0000de",
		16#328f# => X"9ca00001",
		16#3290# => X"a4a500ff",
		16#3291# => X"bc050000",
		16#3292# => X"0c000021",
		16#3293# => X"a88e0001",
		16#3294# => X"a8630001",
		16#3295# => X"e1c27000",
		16#3296# => X"d4022004",
		16#3297# => X"d40e1804",
		16#3298# => X"d4127008",
		16#3299# => X"04000143",
		16#329a# => X"a8700000",
		16#329b# => X"03ffff26",
		16#329c# => X"9d620008",
		16#329d# => X"03ffff59",
		16#329e# => X"9ce7ffff",
		16#329f# => X"e0822000",
		16#32a0# => X"8462000c",
		16#32a1# => X"84a40004",
		16#32a2# => X"84c20008",
		16#32a3# => X"a8a50001",
		16#32a4# => X"d406180c",
		16#32a5# => X"d4033008",
		16#32a6# => X"d4042804",
		16#32a7# => X"04000135",
		16#32a8# => X"a8700000",
		16#32a9# => X"03ffff18",
		16#32aa# => X"9d620008",
		16#32ab# => X"e0822000",
		16#32ac# => X"a8700000",
		16#32ad# => X"84a40004",
		16#32ae# => X"a8a50001",
		16#32af# => X"0400012d",
		16#32b0# => X"d4042804",
		16#32b1# => X"03ffff10",
		16#32b2# => X"9d620008",
		16#32b3# => X"18600001",
		16#32b4# => X"1b800001",
		16#32b5# => X"a863c4bc",
		16#32b6# => X"ab9cb618",
		16#32b7# => X"86c30000",
		16#32b8# => X"847c0000",
		16#32b9# => X"9ed60010",
		16#32ba# => X"bc03ffff",
		16#32bb# => X"10000005",
		16#32bc# => X"e2d67000",
		16#32bd# => X"9ed60fff",
		16#32be# => X"9d60f000",
		16#32bf# => X"e2d65803",
		16#32c0# => X"a8700000",
		16#32c1# => X"040003aa",
		16#32c2# => X"a8960000",
		16#32c3# => X"bc2bffff",
		16#32c4# => X"0c0000ec",
		16#32c5# => X"ab0b0000",
		16#32c6# => X"e082a000",
		16#32c7# => X"e4a45800",
		16#32c8# => X"0c0000a6",
		16#32c9# => X"18a00001",
		16#32ca# => X"1b400001",
		16#32cb# => X"e4245800",
		16#32cc# => X"ab5ac4c8",
		16#32cd# => X"847a0000",
		16#32ce# => X"e0761800",
		16#32cf# => X"0c0000eb",
		16#32d0# => X"d41a1800",
		16#32d1# => X"84bc0000",
		16#32d2# => X"bc25ffff",
		16#32d3# => X"0c0000f9",
		16#32d4# => X"e06b1800",
		16#32d5# => X"e0832002",
		16#32d6# => X"d41a2000",
		16#32d7# => X"a46b0007",
		16#32d8# => X"bc030000",
		16#32d9# => X"10000006",
		16#32da# => X"9c801000",
		16#32db# => X"9c800008",
		16#32dc# => X"e0641802",
		16#32dd# => X"e30b1800",
		16#32de# => X"9c831000",
		16#32df# => X"e2d8b000",
		16#32e0# => X"a8700000",
		16#32e1# => X"a6d60fff",
		16#32e2# => X"e2c4b002",
		16#32e3# => X"04000388",
		16#32e4# => X"a8960000",
		16#32e5# => X"bc0bffff",
		16#32e6# => X"100000e4",
		16#32e7# => X"9c800001",
		16#32e8# => X"e08bc002",
		16#32e9# => X"e084b000",
		16#32ea# => X"a8840001",
		16#32eb# => X"847a0000",
		16#32ec# => X"d4182004",
		16#32ed# => X"e0761800",
		16#32ee# => X"18800001",
		16#32ef# => X"d412c008",
		16#32f0# => X"a884b20c",
		16#32f1# => X"e4022000",
		16#32f2# => X"10000011",
		16#32f3# => X"d41a1800",
		16#32f4# => X"bc54000f",
		16#32f5# => X"0c000099",
		16#32f6# => X"9ca0fff8",
		16#32f7# => X"9c94fff4",
		16#32f8# => X"9cc00005",
		16#32f9# => X"e0842803",
		16#32fa# => X"e0a22000",
		16#32fb# => X"bca4000f",
		16#32fc# => X"d4053004",
		16#32fd# => X"d4053008",
		16#32fe# => X"84a20004",
		16#32ff# => X"a4a50001",
		16#3300# => X"e0842804",
		16#3301# => X"0c0000c2",
		16#3302# => X"d4022004",
		16#3303# => X"18400001",
		16#3304# => X"a842c4c0",
		16#3305# => X"84820000",
		16#3306# => X"e4a32000",
		16#3307# => X"10000003",
		16#3308# => X"18800001",
		16#3309# => X"d4021800",
		16#330a# => X"a884c4c4",
		16#330b# => X"84440000",
		16#330c# => X"e4431000",
		16#330d# => X"0c000065",
		16#330e# => X"15000000",
		16#330f# => X"d4041800",
		16#3310# => X"84520008",
		16#3311# => X"9c60fffc",
		16#3312# => X"84820004",
		16#3313# => X"e0841803",
		16#3314# => X"e0647002",
		16#3315# => X"bda3000f",
		16#3316# => X"10000003",
		16#3317# => X"9ca00001",
		16#3318# => X"9ca00000",
		16#3319# => X"a4a500ff",
		16#331a# => X"bc250000",
		16#331b# => X"10000009",
		16#331c# => X"e44e2000",
		16#331d# => X"10000003",
		16#331e# => X"9cc00001",
		16#331f# => X"a8c50000",
		16#3320# => X"a4c600ff",
		16#3321# => X"bc060000",
		16#3322# => X"13ffff72",
		16#3323# => X"a88e0001",
		16#3324# => X"040000b8",
		16#3325# => X"a8700000",
		16#3326# => X"03fffe9b",
		16#3327# => X"9d600000",
		16#3328# => X"0c00003d",
		16#3329# => X"bc470054",
		16#332a# => X"1000004d",
		16#332b# => X"bc470154",
		16#332c# => X"b8ee004c",
		16#332d# => X"9ce7006e",
		16#332e# => X"03fffeaa",
		16#332f# => X"b8670003",
		16#3330# => X"e0827000",
		16#3331# => X"a9ce0001",
		16#3332# => X"a8e30001",
		16#3333# => X"e0a41800",
		16#3334# => X"d4027004",
		16#3335# => X"d406200c",
		16#3336# => X"d4062008",
		16#3337# => X"d4051800",
		16#3338# => X"d404300c",
		16#3339# => X"d4043008",
		16#333a# => X"d4043804",
		16#333b# => X"040000a1",
		16#333c# => X"a8700000",
		16#333d# => X"03fffe84",
		16#333e# => X"9d620008",
		16#333f# => X"9c620008",
		16#3340# => X"8443000c",
		16#3341# => X"e4031000",
		16#3342# => X"0ffffe71",
		16#3343# => X"9ce70002",
		16#3344# => X"03fffeb4",
		16#3345# => X"18c00001",
		16#3346# => X"e0627000",
		16#3347# => X"84a2000c",
		16#3348# => X"84e20008",
		16#3349# => X"a9ce0001",
		16#334a# => X"d407280c",
		16#334b# => X"d4053808",
		16#334c# => X"e0a32000",
		16#334d# => X"a8e40001",
		16#334e# => X"d406180c",
		16#334f# => X"d4061808",
		16#3350# => X"d4027004",
		16#3351# => X"d403300c",
		16#3352# => X"d4033008",
		16#3353# => X"d4033804",
		16#3354# => X"d4052000",
		16#3355# => X"04000087",
		16#3356# => X"a8700000",
		16#3357# => X"03fffe6a",
		16#3358# => X"9d620008",
		16#3359# => X"e0a22800",
		16#335a# => X"8462000c",
		16#335b# => X"84c50004",
		16#335c# => X"84820008",
		16#335d# => X"a8c60001",
		16#335e# => X"d404180c",
		16#335f# => X"d4032008",
		16#3360# => X"d4053004",
		16#3361# => X"0400007b",
		16#3362# => X"a8700000",
		16#3363# => X"03fffe5e",
		16#3364# => X"9d620008",
		16#3365# => X"9ce7005b",
		16#3366# => X"03fffe72",
		16#3367# => X"b8670003",
		16#3368# => X"10000021",
		16#3369# => X"bc430054",
		16#336a# => X"03fffef7",
		16#336b# => X"9d03005b",
		16#336c# => X"03ffff24",
		16#336d# => X"a8a40000",
		16#336e# => X"a8a5b20c",
		16#336f# => X"e4022800",
		16#3370# => X"13ffff5a",
		16#3371# => X"15000000",
		16#3372# => X"84520008",
		16#3373# => X"9d60fffc",
		16#3374# => X"84820004",
		16#3375# => X"03ffff9f",
		16#3376# => X"e0845803",
		16#3377# => X"1000000c",
		16#3378# => X"bc470554",
		16#3379# => X"b8ee004f",
		16#337a# => X"9ce70077",
		16#337b# => X"03fffe5d",
		16#337c# => X"b8670003",
		16#337d# => X"85720004",
		16#337e# => X"e0a44008",
		16#337f# => X"a8830000",
		16#3380# => X"e0ab2804",
		16#3381# => X"03fffef5",
		16#3382# => X"d4122804",
		16#3383# => X"1000002a",
		16#3384# => X"15000000",
		16#3385# => X"b8ee0052",
		16#3386# => X"9ce7007c",
		16#3387# => X"03fffe51",
		16#3388# => X"b8670003",
		16#3389# => X"1000002c",
		16#338a# => X"bc430154",
		16#338b# => X"b904004c",
		16#338c# => X"03fffed5",
		16#338d# => X"9d08006e",
		16#338e# => X"9c600001",
		16#338f# => X"a8580000",
		16#3390# => X"d4181804",
		16#3391# => X"03ffff83",
		16#3392# => X"9c800000",
		16#3393# => X"a84c0000",
		16#3394# => X"a4a70003",
		16#3395# => X"bc250000",
		16#3396# => X"0c00003f",
		16#3397# => X"9c82fff8",
		16#3398# => X"84420000",
		16#3399# => X"e4222000",
		16#339a# => X"0ffffffa",
		16#339b# => X"9ce7ffff",
		16#339c# => X"e0631800",
		16#339d# => X"84520004",
		16#339e# => X"e4431000",
		16#339f# => X"13fffee2",
		16#33a0# => X"bc030000",
		16#33a1# => X"13fffee0",
		16#33a2# => X"e0831003",
		16#33a3# => X"bc240000",
		16#33a4# => X"13fffe89",
		16#33a5# => X"a8eb0000",
		16#33a6# => X"e0631800",
		16#33a7# => X"e0831003",
		16#33a8# => X"bc040000",
		16#33a9# => X"13fffffd",
		16#33aa# => X"9d6b0004",
		16#33ab# => X"03fffe82",
		16#33ac# => X"a8eb0000",
		16#33ad# => X"9c6003f0",
		16#33ae# => X"03fffe2a",
		16#33af# => X"9ce0007e",
		16#33b0# => X"84520008",
		16#33b1# => X"9c60fffc",
		16#33b2# => X"84820004",
		16#33b3# => X"03ffff61",
		16#33b4# => X"e0841803",
		16#33b5# => X"1000001b",
		16#33b6# => X"bc430554",
		16#33b7# => X"b904004f",
		16#33b8# => X"03fffea9",
		16#33b9# => X"9d080077",
		16#33ba# => X"a4a40fff",
		16#33bb# => X"bc250000",
		16#33bc# => X"13ffff15",
		16#33bd# => X"15000000",
		16#33be# => X"e056a000",
		16#33bf# => X"84920008",
		16#33c0# => X"a8420001",
		16#33c1# => X"03ffff42",
		16#33c2# => X"d4041004",
		16#33c3# => X"9c820008",
		16#33c4# => X"18400001",
		16#33c5# => X"a8700000",
		16#33c6# => X"040016e9",
		16#33c7# => X"a842c4c8",
		16#33c8# => X"03ffff3b",
		16#33c9# => X"84620000",
		16#33ca# => X"03ffff21",
		16#33cb# => X"9ec00000",
		16#33cc# => X"18600001",
		16#33cd# => X"a863b618",
		16#33ce# => X"03ffff09",
		16#33cf# => X"d4035800",
		16#33d0# => X"13fffe91",
		16#33d1# => X"9d00007e",
		16#33d2# => X"b9040052",
		16#33d3# => X"03fffe8e",
		16#33d4# => X"9d08007c",
		16#33d5# => X"84920004",
		16#33d6# => X"ac43ffff",
		16#33d7# => X"e0441003",
		16#33d8# => X"03ffffc4",
		16#33d9# => X"d4121004",
		16#33da# => X"44004800",
		16#33db# => X"15000000",
		16#33dc# => X"44004800",
		16#33dd# => X"15000000",
		16#33de# => X"b4600011",
		16#33df# => X"a8630020",
		16#33e0# => X"c0001840",
		16#33e1# => X"c0004820",
		16#33e2# => X"24000000",
		16#33e3# => X"15000000",
		16#33e4# => X"a8600020",
		16#33e5# => X"ac83ffff",
		16#33e6# => X"b4600011",
		16#33e7# => X"e0641803",
		16#33e8# => X"c0001840",
		16#33e9# => X"c0004820",
		16#33ea# => X"24000000",
		16#33eb# => X"15000000",
		16#33ec# => X"b4600011",
		16#33ed# => X"a8630040",
		16#33ee# => X"c0001840",
		16#33ef# => X"c0004820",
		16#33f0# => X"24000000",
		16#33f1# => X"15000000",
		16#33f2# => X"a8600040",
		16#33f3# => X"ac83ffff",
		16#33f4# => X"b4600011",
		16#33f5# => X"e0641803",
		16#33f6# => X"c0001840",
		16#33f7# => X"c0004820",
		16#33f8# => X"24000000",
		16#33f9# => X"15000000",
		16#33fa# => X"b4600001",
		16#33fb# => X"a4830004",
		16#33fc# => X"e4040000",
		16#33fd# => X"10000021",
		16#33fe# => X"15000000",
		16#33ff# => X"b4c00011",
		16#3400# => X"9ca0ffff",
		16#3401# => X"aca50010",
		16#3402# => X"e0a62803",
		16#3403# => X"c0002811",
		16#3404# => X"b4600006",
		16#3405# => X"a4830080",
		16#3406# => X"b8e40047",
		16#3407# => X"a9000010",
		16#3408# => X"e1c83808",
		16#3409# => X"a4830078",
		16#340a# => X"b8e40043",
		16#340b# => X"a9000001",
		16#340c# => X"e1a83808",
		16#340d# => X"9cc00000",
		16#340e# => X"e0ae3808",
		16#340f# => X"c0803002",
		16#3410# => X"e4262800",
		16#3411# => X"13fffffe",
		16#3412# => X"e0c67000",
		16#3413# => X"b4c00011",
		16#3414# => X"a8c60010",
		16#3415# => X"c0003011",
		16#3416# => X"15000000",
		16#3417# => X"15000000",
		16#3418# => X"15000000",
		16#3419# => X"15000000",
		16#341a# => X"15000000",
		16#341b# => X"15000000",
		16#341c# => X"15000000",
		16#341d# => X"15000000",
		16#341e# => X"b4600001",
		16#341f# => X"a4830002",
		16#3420# => X"e4040000",
		16#3421# => X"10000019",
		16#3422# => X"15000000",
		16#3423# => X"b4c00011",
		16#3424# => X"9ca0ffff",
		16#3425# => X"aca50008",
		16#3426# => X"e0a62803",
		16#3427# => X"c0002811",
		16#3428# => X"b4600005",
		16#3429# => X"a4830080",
		16#342a# => X"b8e40047",
		16#342b# => X"a9000010",
		16#342c# => X"e1c83808",
		16#342d# => X"a4830078",
		16#342e# => X"b8e40043",
		16#342f# => X"a9000001",
		16#3430# => X"e1a83808",
		16#3431# => X"9cc00000",
		16#3432# => X"e0ae3808",
		16#3433# => X"c0603003",
		16#3434# => X"e4262800",
		16#3435# => X"13fffffe",
		16#3436# => X"e0c67000",
		16#3437# => X"b4c00011",
		16#3438# => X"a8c60008",
		16#3439# => X"c0003011",
		16#343a# => X"44004800",
		16#343b# => X"15000000",
		16#343c# => X"b5a00011",
		16#343d# => X"a9ad0010",
		16#343e# => X"c0006811",
		16#343f# => X"15000000",
		16#3440# => X"15000000",
		16#3441# => X"15000000",
		16#3442# => X"15000000",
		16#3443# => X"15000000",
		16#3444# => X"44004800",
		16#3445# => X"15000000",
		16#3446# => X"b5a00011",
		16#3447# => X"9d80ffff",
		16#3448# => X"ad8c0010",
		16#3449# => X"e18d6003",
		16#344a# => X"c0006011",
		16#344b# => X"44004800",
		16#344c# => X"15000000",
		16#344d# => X"44004800",
		16#344e# => X"c0801802",
		16#344f# => X"b5a00011",
		16#3450# => X"a9ad0008",
		16#3451# => X"c0006811",
		16#3452# => X"15000000",
		16#3453# => X"15000000",
		16#3454# => X"15000000",
		16#3455# => X"15000000",
		16#3456# => X"15000000",
		16#3457# => X"44004800",
		16#3458# => X"15000000",
		16#3459# => X"b5a00011",
		16#345a# => X"9d80ffff",
		16#345b# => X"ad8c0008",
		16#345c# => X"e18d6003",
		16#345d# => X"c0006011",
		16#345e# => X"44004800",
		16#345f# => X"15000000",
		16#3460# => X"44004800",
		16#3461# => X"c0601803",
		16#3462# => X"9c21fff4",
		16#3463# => X"d4014800",
		16#3464# => X"b4604802",
		16#3465# => X"18e00001",
		16#3466# => X"a8e7b61c",
		16#3467# => X"1900ffff",
		16#3468# => X"a908ffff",
		16#3469# => X"19800001",
		16#346a# => X"a98cb69c",
		16#346b# => X"e083000f",
		16#346c# => X"e4240000",
		16#346d# => X"0c000014",
		16#346e# => X"15000000",
		16#346f# => X"9ca4ffff",
		16#3470# => X"b8c50002",
		16#3471# => X"e1c63800",
		16#3472# => X"e1a66000",
		16#3473# => X"85ce0000",
		16#3474# => X"e42e4000",
		16#3475# => X"0c000008",
		16#3476# => X"15000000",
		16#3477# => X"d4011804",
		16#3478# => X"846d0000",
		16#3479# => X"48007000",
		16#347a# => X"d4012808",
		16#347b# => X"84610004",
		16#347c# => X"84a10008",
		16#347d# => X"a8c00001",
		16#347e# => X"e0c62808",
		16#347f# => X"03ffffec",
		16#3480# => X"e0633005",
		16#3481# => X"85210000",
		16#3482# => X"c1201802",
		16#3483# => X"44004800",
		16#3484# => X"9c21000c",
		16#3485# => X"9c21fffc",
		16#3486# => X"d4013000",
		16#3487# => X"b8630002",
		16#3488# => X"18c00001",
		16#3489# => X"a8c6b61c",
		16#348a# => X"e0c61800",
		16#348b# => X"d4062000",
		16#348c# => X"18c00001",
		16#348d# => X"a8c6b69c",
		16#348e# => X"e0c61800",
		16#348f# => X"d4062800",
		16#3490# => X"84c10000",
		16#3491# => X"44004800",
		16#3492# => X"9c210004",
		16#3493# => X"9c21fffc",
		16#3494# => X"d4012000",
		16#3495# => X"a8800001",
		16#3496# => X"e0841808",
		16#3497# => X"b4604800",
		16#3498# => X"e0632004",
		16#3499# => X"c1201800",
		16#349a# => X"84810000",
		16#349b# => X"44004800",
		16#349c# => X"9c210004",
		16#349d# => X"9c21fffc",
		16#349e# => X"d4012000",
		16#349f# => X"a8800001",
		16#34a0# => X"e0841808",
		16#34a1# => X"ac84ffff",
		16#34a2# => X"b4604800",
		16#34a3# => X"e0632003",
		16#34a4# => X"c1201800",
		16#34a5# => X"84810000",
		16#34a6# => X"44004800",
		16#34a7# => X"9c210004",
		16#34a8# => X"d4011000",
		16#34a9# => X"d401280c",
		16#34aa# => X"d4013010",
		16#34ab# => X"d4013814",
		16#34ac# => X"d4014018",
		16#34ad# => X"d401481c",
		16#34ae# => X"d4015020",
		16#34af# => X"d4015824",
		16#34b0# => X"d4016028",
		16#34b1# => X"d401682c",
		16#34b2# => X"d4017030",
		16#34b3# => X"d4017834",
		16#34b4# => X"d4018038",
		16#34b5# => X"d401883c",
		16#34b6# => X"d4019040",
		16#34b7# => X"d4019844",
		16#34b8# => X"d401a048",
		16#34b9# => X"d401a84c",
		16#34ba# => X"d401b050",
		16#34bb# => X"d401b854",
		16#34bc# => X"d401c058",
		16#34bd# => X"d401c85c",
		16#34be# => X"d401d060",
		16#34bf# => X"d401d864",
		16#34c0# => X"d401e068",
		16#34c1# => X"d401e86c",
		16#34c2# => X"d401f070",
		16#34c3# => X"d401f874",
		16#34c4# => X"a5a3ffff",
		16#34c5# => X"b9ad0046",
		16#34c6# => X"9dadfff8",
		16#34c7# => X"19c00001",
		16#34c8# => X"a9ceb71c",
		16#34c9# => X"e1ce6800",
		16#34ca# => X"85ae0000",
		16#34cb# => X"19e0ffff",
		16#34cc# => X"a9efffff",
		16#34cd# => X"e42d7800",
		16#34ce# => X"0c000025",
		16#34cf# => X"15000000",
		16#34d0# => X"48006800",
		16#34d1# => X"e0642004",
		16#34d2# => X"84410000",
		16#34d3# => X"84610004",
		16#34d4# => X"84810008",
		16#34d5# => X"84a1000c",
		16#34d6# => X"84c10010",
		16#34d7# => X"84e10014",
		16#34d8# => X"85010018",
		16#34d9# => X"8521001c",
		16#34da# => X"85410020",
		16#34db# => X"85610024",
		16#34dc# => X"85810028",
		16#34dd# => X"85a1002c",
		16#34de# => X"85c10030",
		16#34df# => X"85e10034",
		16#34e0# => X"86010038",
		16#34e1# => X"8621003c",
		16#34e2# => X"86410040",
		16#34e3# => X"86610044",
		16#34e4# => X"86810048",
		16#34e5# => X"86a1004c",
		16#34e6# => X"86c10050",
		16#34e7# => X"86e10054",
		16#34e8# => X"87010058",
		16#34e9# => X"8721005c",
		16#34ea# => X"87410060",
		16#34eb# => X"87610064",
		16#34ec# => X"87810068",
		16#34ed# => X"87a1006c",
		16#34ee# => X"87c10070",
		16#34ef# => X"87e10074",
		16#34f0# => X"9c210100",
		16#34f1# => X"24000000",
		16#34f2# => X"15000000",
		16#34f3# => X"07fffc72",
		16#34f4# => X"e0642004",
		16#34f5# => X"9c21fffc",
		16#34f6# => X"d4012800",
		16#34f7# => X"b8630002",
		16#34f8# => X"9c63fff8",
		16#34f9# => X"18a00001",
		16#34fa# => X"a8a5b71c",
		16#34fb# => X"e0a51800",
		16#34fc# => X"d4052000",
		16#34fd# => X"84a10000",
		16#34fe# => X"44004800",
		16#34ff# => X"9c210004",
		16#3500# => X"18600001",
		16#3501# => X"18800001",
		16#3502# => X"a863c500",
		16#3503# => X"d7e117fc",
		16#3504# => X"a884c504",
		16#3505# => X"18400fff",
		16#3506# => X"84a30000",
		16#3507# => X"84840000",
		16#3508# => X"a842ffff",
		16#3509# => X"9ca50001",
		16#350a# => X"e0841003",
		16#350b# => X"18406000",
		16#350c# => X"d4032800",
		16#350d# => X"9c21fffc",
		16#350e# => X"e0841004",
		16#350f# => X"9c605000",
		16#3510# => X"c0032000",
		16#3511# => X"9c210004",
		16#3512# => X"44004800",
		16#3513# => X"8441fffc",
		16#3514# => X"9c630000",
		16#3515# => X"15000002",
		16#3516# => X"44004800",
		16#3517# => X"15000000",
		16#3518# => X"c0032000",
		16#3519# => X"44004800",
		16#351a# => X"15000000",
		16#351b# => X"b5630000",
		16#351c# => X"44004800",
		16#351d# => X"15000000",
		16#351e# => X"18600001",
		16#351f# => X"d7e117fc",
		16#3520# => X"a863b790",
		16#3521# => X"18800001",
		16#3522# => X"84a30000",
		16#3523# => X"1840d000",
		16#3524# => X"a5650001",
		16#3525# => X"a884c4f0",
		16#3526# => X"a8420001",
		16#3527# => X"e1605802",
		16#3528# => X"b8a50041",
		16#3529# => X"84c40000",
		16#352a# => X"e16b1003",
		16#352b# => X"9cc60001",
		16#352c# => X"e16b2805",
		16#352d# => X"9c21fffc",
		16#352e# => X"d4043000",
		16#352f# => X"d4035800",
		16#3530# => X"9c210004",
		16#3531# => X"44004800",
		16#3532# => X"8441fffc",
		16#3533# => X"a8830000",
		16#3534# => X"18600001",
		16#3535# => X"d7e14ffc",
		16#3536# => X"a8637da4",
		16#3537# => X"d7e117f8",
		16#3538# => X"84630000",
		16#3539# => X"9c21fff8",
		16#353a# => X"07fff092",
		16#353b# => X"9c400000",
		16#353c# => X"18a00001",
		16#353d# => X"18800000",
		16#353e# => X"a8a5c504",
		16#353f# => X"9c600005",
		16#3540# => X"d4055800",
		16#3541# => X"18a00001",
		16#3542# => X"a884d400",
		16#3543# => X"a8a5c500",
		16#3544# => X"d4051000",
		16#3545# => X"9c210008",
		16#3546# => X"8521fffc",
		16#3547# => X"03ffffae",
		16#3548# => X"8441fff8",
		16#3549# => X"18600001",
		16#354a# => X"d7e117fc",
		16#354b# => X"a863c504",
		16#354c# => X"18400fff",
		16#354d# => X"84830000",
		16#354e# => X"a842ffff",
		16#354f# => X"9c21fffc",
		16#3550# => X"e0841003",
		16#3551# => X"18406000",
		16#3552# => X"9c605000",
		16#3553# => X"e0841004",
		16#3554# => X"c0032000",
		16#3555# => X"9c600011",
		16#3556# => X"b4830000",
		16#3557# => X"a8840002",
		16#3558# => X"c0032000",
		16#3559# => X"9c210004",
		16#355a# => X"44004800",
		16#355b# => X"8441fffc",
		16#355c# => X"d7e117fc",
		16#355d# => X"9c600011",
		16#355e# => X"9c21fffc",
		16#355f# => X"b4830000",
		16#3560# => X"9c40fffd",
		16#3561# => X"e0841003",
		16#3562# => X"c0032000",
		16#3563# => X"9c210004",
		16#3564# => X"44004800",
		16#3565# => X"8441fffc",
		16#3566# => X"18600001",
		16#3567# => X"a863c500",
		16#3568# => X"85630000",
		16#3569# => X"44004800",
		16#356a# => X"15000000",
		16#356b# => X"18600001",
		16#356c# => X"d7e117fc",
		16#356d# => X"a863c500",
		16#356e# => X"9c400000",
		16#356f# => X"9c21fffc",
		16#3570# => X"d4031000",
		16#3571# => X"9c210004",
		16#3572# => X"44004800",
		16#3573# => X"8441fffc",
		16#3574# => X"d7e14ffc",
		16#3575# => X"9c21fffc",
		16#3576# => X"a8a40000",
		16#3577# => X"9cc10004",
		16#3578# => X"0400014e",
		16#3579# => X"84830008",
		16#357a# => X"9c210004",
		16#357b# => X"8521fffc",
		16#357c# => X"44004800",
		16#357d# => X"15000000",
		16#357e# => X"a8a30000",
		16#357f# => X"18600001",
		16#3580# => X"d7e14ffc",
		16#3581# => X"a863ade4",
		16#3582# => X"9c21fffc",
		16#3583# => X"84630000",
		16#3584# => X"9cc10004",
		16#3585# => X"04000141",
		16#3586# => X"84830008",
		16#3587# => X"9c210004",
		16#3588# => X"8521fffc",
		16#3589# => X"44004800",
		16#358a# => X"15000000",
		16#358b# => X"d7e14ffc",
		16#358c# => X"9c21fffc",
		16#358d# => X"84a30008",
		16#358e# => X"9c210004",
		16#358f# => X"8521fffc",
		16#3590# => X"0000000d",
		16#3591# => X"15000000",
		16#3592# => X"a8830000",
		16#3593# => X"18600001",
		16#3594# => X"d7e14ffc",
		16#3595# => X"a863ade4",
		16#3596# => X"9c21fffc",
		16#3597# => X"84630000",
		16#3598# => X"84a30008",
		16#3599# => X"9c210004",
		16#359a# => X"8521fffc",
		16#359b# => X"00000002",
		16#359c# => X"15000000",
		16#359d# => X"d7e117f0",
		16#359e# => X"d7e177f4",
		16#359f# => X"d7e187f8",
		16#35a0# => X"d7e14ffc",
		16#35a1# => X"a9c30000",
		16#35a2# => X"9c21fff0",
		16#35a3# => X"aa040000",
		16#35a4# => X"bc030000",
		16#35a5# => X"10000006",
		16#35a6# => X"a8450000",
		16#35a7# => X"84830038",
		16#35a8# => X"bc240000",
		16#35a9# => X"0c000026",
		16#35aa# => X"15000000",
		16#35ab# => X"84620008",
		16#35ac# => X"9c63ffff",
		16#35ad# => X"bd630000",
		16#35ae# => X"0c00000e",
		16#35af# => X"d4021808",
		16#35b0# => X"84620000",
		16#35b1# => X"d8038000",
		16#35b2# => X"84820000",
		16#35b3# => X"9c640001",
		16#35b4# => X"8d640000",
		16#35b5# => X"d4021800",
		16#35b6# => X"9c210010",
		16#35b7# => X"8521fffc",
		16#35b8# => X"8441fff0",
		16#35b9# => X"85c1fff4",
		16#35ba# => X"44004800",
		16#35bb# => X"8601fff8",
		16#35bc# => X"84820018",
		16#35bd# => X"e5832000",
		16#35be# => X"10000015",
		16#35bf# => X"a86e0000",
		16#35c0# => X"84620000",
		16#35c1# => X"d8038000",
		16#35c2# => X"84620000",
		16#35c3# => X"8c830000",
		16#35c4# => X"bc04000a",
		16#35c5# => X"10000016",
		16#35c6# => X"9c630001",
		16#35c7# => X"a9640000",
		16#35c8# => X"d4021800",
		16#35c9# => X"9c210010",
		16#35ca# => X"8521fffc",
		16#35cb# => X"8441fff0",
		16#35cc# => X"85c1fff4",
		16#35cd# => X"44004800",
		16#35ce# => X"8601fff8",
		16#35cf# => X"040013bf",
		16#35d0# => X"15000000",
		16#35d1# => X"03ffffdb",
		16#35d2# => X"84620008",
		16#35d3# => X"9c210010",
		16#35d4# => X"a8900000",
		16#35d5# => X"a8a20000",
		16#35d6# => X"8521fffc",
		16#35d7# => X"8441fff0",
		16#35d8# => X"85c1fff4",
		16#35d9# => X"00000938",
		16#35da# => X"8601fff8",
		16#35db# => X"9c210010",
		16#35dc# => X"a86e0000",
		16#35dd# => X"a8a20000",
		16#35de# => X"8521fffc",
		16#35df# => X"8441fff0",
		16#35e0# => X"85c1fff4",
		16#35e1# => X"00000930",
		16#35e2# => X"8601fff8",
		16#35e3# => X"d7e187f8",
		16#35e4# => X"1a000001",
		16#35e5# => X"d7e117f0",
		16#35e6# => X"aa10ade4",
		16#35e7# => X"d7e177f4",
		16#35e8# => X"d7e14ffc",
		16#35e9# => X"84b00000",
		16#35ea# => X"9c21fff0",
		16#35eb# => X"a9c30000",
		16#35ec# => X"bc050000",
		16#35ed# => X"10000006",
		16#35ee# => X"a8440000",
		16#35ef# => X"84650038",
		16#35f0# => X"bc230000",
		16#35f1# => X"0c000026",
		16#35f2# => X"15000000",
		16#35f3# => X"84620008",
		16#35f4# => X"9c63ffff",
		16#35f5# => X"bd630000",
		16#35f6# => X"0c00000e",
		16#35f7# => X"d4021808",
		16#35f8# => X"84620000",
		16#35f9# => X"d8037000",
		16#35fa# => X"84820000",
		16#35fb# => X"9c640001",
		16#35fc# => X"8d640000",
		16#35fd# => X"d4021800",
		16#35fe# => X"9c210010",
		16#35ff# => X"8521fffc",
		16#3600# => X"8441fff0",
		16#3601# => X"85c1fff4",
		16#3602# => X"44004800",
		16#3603# => X"8601fff8",
		16#3604# => X"84820018",
		16#3605# => X"e5832000",
		16#3606# => X"10000015",
		16#3607# => X"a88e0000",
		16#3608# => X"84620000",
		16#3609# => X"d8037000",
		16#360a# => X"84620000",
		16#360b# => X"8c830000",
		16#360c# => X"bc04000a",
		16#360d# => X"10000016",
		16#360e# => X"9c630001",
		16#360f# => X"a9640000",
		16#3610# => X"d4021800",
		16#3611# => X"9c210010",
		16#3612# => X"8521fffc",
		16#3613# => X"8441fff0",
		16#3614# => X"85c1fff4",
		16#3615# => X"44004800",
		16#3616# => X"8601fff8",
		16#3617# => X"04001377",
		16#3618# => X"a8650000",
		16#3619# => X"03ffffdb",
		16#361a# => X"84620008",
		16#361b# => X"84700000",
		16#361c# => X"9c210010",
		16#361d# => X"a8a20000",
		16#361e# => X"8521fffc",
		16#361f# => X"8441fff0",
		16#3620# => X"85c1fff4",
		16#3621# => X"000008f0",
		16#3622# => X"8601fff8",
		16#3623# => X"84700000",
		16#3624# => X"9c210010",
		16#3625# => X"a8a20000",
		16#3626# => X"8521fffc",
		16#3627# => X"8441fff0",
		16#3628# => X"85c1fff4",
		16#3629# => X"000008e8",
		16#362a# => X"8601fff8",
		16#362b# => X"d7e117f4",
		16#362c# => X"d7e177f8",
		16#362d# => X"d7e14ffc",
		16#362e# => X"a8430000",
		16#362f# => X"9c21ffd8",
		16#3630# => X"a8640000",
		16#3631# => X"04000057",
		16#3632# => X"a9c40000",
		16#3633# => X"18600001",
		16#3634# => X"18e00001",
		16#3635# => X"a863ade4",
		16#3636# => X"9ccb0001",
		16#3637# => X"84630000",
		16#3638# => X"a8e7853a",
		16#3639# => X"84a30008",
		16#363a# => X"d4013808",
		16#363b# => X"9865000c",
		16#363c# => X"9ce00001",
		16#363d# => X"d4013018",
		16#363e# => X"9cc00002",
		16#363f# => X"a4832000",
		16#3640# => X"d4017000",
		16#3641# => X"d4015804",
		16#3642# => X"d401380c",
		16#3643# => X"d4010810",
		16#3644# => X"bc240000",
		16#3645# => X"10000008",
		16#3646# => X"d4013014",
		16#3647# => X"84850064",
		16#3648# => X"9cc0dfff",
		16#3649# => X"a8632000",
		16#364a# => X"e0843003",
		16#364b# => X"dc05180c",
		16#364c# => X"d4052064",
		16#364d# => X"a8620000",
		16#364e# => X"9ca10010",
		16#364f# => X"0400152c",
		16#3650# => X"84820008",
		16#3651# => X"bc0b0000",
		16#3652# => X"0c000008",
		16#3653# => X"9c60000a",
		16#3654# => X"9c210028",
		16#3655# => X"a9630000",
		16#3656# => X"8521fffc",
		16#3657# => X"8441fff4",
		16#3658# => X"44004800",
		16#3659# => X"85c1fff8",
		16#365a# => X"9c210028",
		16#365b# => X"9c60ffff",
		16#365c# => X"8521fffc",
		16#365d# => X"a9630000",
		16#365e# => X"8441fff4",
		16#365f# => X"44004800",
		16#3660# => X"85c1fff8",
		16#3661# => X"a8830000",
		16#3662# => X"18600001",
		16#3663# => X"d7e14ffc",
		16#3664# => X"a863ade4",
		16#3665# => X"9c21fffc",
		16#3666# => X"84630000",
		16#3667# => X"9c210004",
		16#3668# => X"8521fffc",
		16#3669# => X"03ffffc2",
		16#366a# => X"15000000",
		16#366b# => X"d7e117f4",
		16#366c# => X"18400001",
		16#366d# => X"d7e177f8",
		16#366e# => X"a842c508",
		16#366f# => X"a9c30000",
		16#3670# => X"a8640000",
		16#3671# => X"9c800000",
		16#3672# => X"d7e14ffc",
		16#3673# => X"d4022000",
		16#3674# => X"04002853",
		16#3675# => X"9c21fff4",
		16#3676# => X"bc2bffff",
		16#3677# => X"0c000007",
		16#3678# => X"15000000",
		16#3679# => X"9c21000c",
		16#367a# => X"8521fffc",
		16#367b# => X"8441fff4",
		16#367c# => X"44004800",
		16#367d# => X"85c1fff8",
		16#367e# => X"84420000",
		16#367f# => X"bc020000",
		16#3680# => X"13fffff9",
		16#3681# => X"15000000",
		16#3682# => X"d40e1000",
		16#3683# => X"9c21000c",
		16#3684# => X"8521fffc",
		16#3685# => X"8441fff4",
		16#3686# => X"44004800",
		16#3687# => X"85c1fff8",
		16#3688# => X"d7e117fc",
		16#3689# => X"a4830003",
		16#368a# => X"bc040000",
		16#368b# => X"10000039",
		16#368c# => X"9c21fffc",
		16#368d# => X"91630000",
		16#368e# => X"bc0b0000",
		16#368f# => X"10000032",
		16#3690# => X"15000000",
		16#3691# => X"00000006",
		16#3692# => X"a9630000",
		16#3693# => X"908b0000",
		16#3694# => X"bc240000",
		16#3695# => X"0c00002b",
		16#3696# => X"15000000",
		16#3697# => X"9d6b0001",
		16#3698# => X"a48b0003",
		16#3699# => X"bc240000",
		16#369a# => X"13fffff9",
		16#369b# => X"15000000",
		16#369c# => X"1840fefe",
		16#369d# => X"848b0000",
		16#369e# => X"a842feff",
		16#369f# => X"e0a41000",
		16#36a0# => X"ac84ffff",
		16#36a1# => X"18408080",
		16#36a2# => X"e0852003",
		16#36a3# => X"a8428080",
		16#36a4# => X"e0841003",
		16#36a5# => X"bc240000",
		16#36a6# => X"10000010",
		16#36a7# => X"15000000",
		16#36a8# => X"9d6b0004",
		16#36a9# => X"1840fefe",
		16#36aa# => X"848b0000",
		16#36ab# => X"a842feff",
		16#36ac# => X"e0a41000",
		16#36ad# => X"ac84ffff",
		16#36ae# => X"18408080",
		16#36af# => X"e0852003",
		16#36b0# => X"a8428080",
		16#36b1# => X"e0841003",
		16#36b2# => X"bc040000",
		16#36b3# => X"13fffff6",
		16#36b4# => X"9d6b0004",
		16#36b5# => X"9d6bfffc",
		16#36b6# => X"908b0000",
		16#36b7# => X"bc040000",
		16#36b8# => X"10000008",
		16#36b9# => X"15000000",
		16#36ba# => X"9d6b0001",
		16#36bb# => X"908b0000",
		16#36bc# => X"bc240000",
		16#36bd# => X"13fffffe",
		16#36be# => X"9d6b0001",
		16#36bf# => X"9d6bffff",
		16#36c0# => X"e16b1802",
		16#36c1# => X"9c210004",
		16#36c2# => X"44004800",
		16#36c3# => X"8441fffc",
		16#36c4# => X"03ffffd8",
		16#36c5# => X"a9630000",
		16#36c6# => X"d7e14ffc",
		16#36c7# => X"d7e117d4",
		16#36c8# => X"d7e177d8",
		16#36c9# => X"d7e187dc",
		16#36ca# => X"d7e197e0",
		16#36cb# => X"d7e1a7e4",
		16#36cc# => X"d7e1b7e8",
		16#36cd# => X"d7e1c7ec",
		16#36ce# => X"d7e1d7f0",
		16#36cf# => X"d7e1e7f4",
		16#36d0# => X"d7e1f7f8",
		16#36d1# => X"9c21fa78",
		16#36d2# => X"a9c50000",
		16#36d3# => X"d4011828",
		16#36d4# => X"d4012020",
		16#36d5# => X"040016ab",
		16#36d6# => X"d401302c",
		16#36d7# => X"856b0000",
		16#36d8# => X"a86b0000",
		16#36d9# => X"07ffffaf",
		16#36da# => X"d4015848",
		16#36db# => X"84410028",
		16#36dc# => X"bc020000",
		16#36dd# => X"10000006",
		16#36de# => X"d4015854",
		16#36df# => X"84420038",
		16#36e0# => X"bc220000",
		16#36e1# => X"0c00012d",
		16#36e2# => X"15000000",
		16#36e3# => X"84610020",
		16#36e4# => X"9843000c",
		16#36e5# => X"a4e2ffff",
		16#36e6# => X"a4a72000",
		16#36e7# => X"bc250000",
		16#36e8# => X"1000000b",
		16#36e9# => X"a4a70008",
		16#36ea# => X"84a30064",
		16#36eb# => X"9c60dfff",
		16#36ec# => X"a8422000",
		16#36ed# => X"84810020",
		16#36ee# => X"e0a51803",
		16#36ef# => X"dc04100c",
		16#36f0# => X"d4042864",
		16#36f1# => X"a4e2ffff",
		16#36f2# => X"a4a70008",
		16#36f3# => X"bc050000",
		16#36f4# => X"1000076f",
		16#36f5# => X"84810020",
		16#36f6# => X"84a40010",
		16#36f7# => X"bc250000",
		16#36f8# => X"0c00076c",
		16#36f9# => X"84610028",
		16#36fa# => X"a4e7001a",
		16#36fb# => X"bc27000a",
		16#36fc# => X"0c0000e5",
		16#36fd# => X"84610020",
		16#36fe# => X"9c400000",
		16#36ff# => X"9c610538",
		16#3700# => X"9c810537",
		16#3701# => X"d4011814",
		16#3702# => X"d4012010",
		16#3703# => X"9c600000",
		16#3704# => X"d4011038",
		16#3705# => X"9c4104d0",
		16#3706# => X"d4011d40",
		16#3707# => X"d4011538",
		16#3708# => X"d4011d3c",
		16#3709# => X"d401184c",
		16#370a# => X"d4011850",
		16#370b# => X"d401185c",
		16#370c# => X"d4011858",
		16#370d# => X"d4011830",
		16#370e# => X"aac20000",
		16#370f# => X"84610010",
		16#3710# => X"84410014",
		16#3711# => X"9c810544",
		16#3712# => X"e0421802",
		16#3713# => X"d401701c",
		16#3714# => X"d4011064",
		16#3715# => X"9c41046f",
		16#3716# => X"d4012008",
		16#3717# => X"d401100c",
		16#3718# => X"8461001c",
		16#3719# => X"90a30000",
		16#371a# => X"ac450025",
		16#371b# => X"a44200ff",
		16#371c# => X"bc020000",
		16#371d# => X"100000f5",
		16#371e# => X"a44500ff",
		16#371f# => X"bc020000",
		16#3720# => X"100000f2",
		16#3721# => X"15000000",
		16#3722# => X"00000005",
		16#3723# => X"a9c30000",
		16#3724# => X"bc220000",
		16#3725# => X"0c00000a",
		16#3726# => X"8481001c",
		16#3727# => X"9dce0001",
		16#3728# => X"90ae0000",
		16#3729# => X"ac450025",
		16#372a# => X"a44200ff",
		16#372b# => X"bc020000",
		16#372c# => X"0ffffff8",
		16#372d# => X"a44500ff",
		16#372e# => X"8481001c",
		16#372f# => X"e04e2002",
		16#3730# => X"bc020000",
		16#3731# => X"10000010",
		16#3732# => X"86410540",
		16#3733# => X"8601053c",
		16#3734# => X"e2521000",
		16#3735# => X"9e100001",
		16#3736# => X"d4162000",
		16#3737# => X"d4161004",
		16#3738# => X"d4019540",
		16#3739# => X"bd500007",
		16#373a# => X"10000080",
		16#373b# => X"d401853c",
		16#373c# => X"9ed60008",
		16#373d# => X"84610030",
		16#373e# => X"e0631000",
		16#373f# => X"d4011830",
		16#3740# => X"90ae0000",
		16#3741# => X"bc050000",
		16#3742# => X"10000081",
		16#3743# => X"9d000000",
		16#3744# => X"9dce0001",
		16#3745# => X"9c800000",
		16#3746# => X"d401701c",
		16#3747# => X"d801255b",
		16#3748# => X"9e40ffff",
		16#3749# => X"d4014034",
		16#374a# => X"d4014018",
		16#374b# => X"a8ae0000",
		16#374c# => X"93c50000",
		16#374d# => X"9ca50001",
		16#374e# => X"9c7effe0",
		16#374f# => X"bc430058",
		16#3750# => X"0c000056",
		16#3751# => X"18400001",
		16#3752# => X"d401281c",
		16#3753# => X"bc1e0000",
		16#3754# => X"1000006f",
		16#3755# => X"d801455b",
		16#3756# => X"9c800001",
		16#3757# => X"9c400000",
		16#3758# => X"9c610510",
		16#3759# => X"d4012024",
		16#375a# => X"d801f510",
		16#375b# => X"d801155b",
		16#375c# => X"ab440000",
		16#375d# => X"d4011840",
		16#375e# => X"9c400000",
		16#375f# => X"d4011044",
		16#3760# => X"84410018",
		16#3761# => X"a7820002",
		16#3762# => X"bc1c0000",
		16#3763# => X"10000006",
		16#3764# => X"84810018",
		16#3765# => X"84610024",
		16#3766# => X"9c630002",
		16#3767# => X"d4011824",
		16#3768# => X"84810018",
		16#3769# => X"a4840084",
		16#376a# => X"bc040000",
		16#376b# => X"0c00022a",
		16#376c# => X"d401203c",
		16#376d# => X"84410034",
		16#376e# => X"84610024",
		16#376f# => X"e1c21802",
		16#3770# => X"bd4e0000",
		16#3771# => X"0c000224",
		16#3772# => X"bd4e0010",
		16#3773# => X"0c0006ce",
		16#3774# => X"15000000",
		16#3775# => X"1a800001",
		16#3776# => X"d401e060",
		16#3777# => X"86410540",
		16#3778# => X"ab9a0000",
		16#3779# => X"8601053c",
		16#377a# => X"aa948a4c",
		16#377b# => X"9f000010",
		16#377c# => X"84410028",
		16#377d# => X"00000007",
		16#377e# => X"87410020",
		16#377f# => X"9ed60008",
		16#3780# => X"9dcefff0",
		16#3781# => X"bd4e0010",
		16#3782# => X"0c000017",
		16#3783# => X"9cf60008",
		16#3784# => X"9e100001",
		16#3785# => X"9e520010",
		16#3786# => X"d416a000",
		16#3787# => X"d416c004",
		16#3788# => X"d4019540",
		16#3789# => X"bd500007",
		16#378a# => X"0ffffff5",
		16#378b# => X"d401853c",
		16#378c# => X"a8620000",
		16#378d# => X"a89a0000",
		16#378e# => X"04001f88",
		16#378f# => X"9ca10538",
		16#3790# => X"bc2b0000",
		16#3791# => X"1000003a",
		16#3792# => X"9dcefff0",
		16#3793# => X"9ce104d8",
		16#3794# => X"9ec104d0",
		16#3795# => X"86410540",
		16#3796# => X"bd4e0010",
		16#3797# => X"13ffffed",
		16#3798# => X"8601053c",
		16#3799# => X"ab5c0000",
		16#379a# => X"87810060",
		16#379b# => X"9e100001",
		16#379c# => X"e2527000",
		16#379d# => X"d416a000",
		16#379e# => X"d4167004",
		16#379f# => X"d4019540",
		16#37a0# => X"bd500007",
		16#37a1# => X"10000447",
		16#37a2# => X"d401853c",
		16#37a3# => X"9f070008",
		16#37a4# => X"000001f4",
		16#37a5# => X"aac70000",
		16#37a6# => X"b8630002",
		16#37a7# => X"a84288d8",
		16#37a8# => X"e0631000",
		16#37a9# => X"84630000",
		16#37aa# => X"44001800",
		16#37ab# => X"15000000",
		16#37ac# => X"8441002c",
		16#37ad# => X"8461002c",
		16#37ae# => X"84420000",
		16#37af# => X"9c630004",
		16#37b0# => X"d4011034",
		16#37b1# => X"bd620000",
		16#37b2# => X"13ffff9a",
		16#37b3# => X"d401182c",
		16#37b4# => X"e0401002",
		16#37b5# => X"d4011034",
		16#37b6# => X"84810018",
		16#37b7# => X"a8840004",
		16#37b8# => X"03ffff94",
		16#37b9# => X"d4012018",
		16#37ba# => X"84610028",
		16#37bb# => X"84810020",
		16#37bc# => X"04001f5a",
		16#37bd# => X"9ca10538",
		16#37be# => X"bc2b0000",
		16#37bf# => X"1000000c",
		16#37c0# => X"9ec104d0",
		16#37c1# => X"03ffff7d",
		16#37c2# => X"84610030",
		16#37c3# => X"84410540",
		16#37c4# => X"bc020000",
		16#37c5# => X"10000007",
		16#37c6# => X"84610020",
		16#37c7# => X"84610028",
		16#37c8# => X"84810020",
		16#37c9# => X"04001f4d",
		16#37ca# => X"9ca10538",
		16#37cb# => X"84610020",
		16#37cc# => X"9443000c",
		16#37cd# => X"a4420040",
		16#37ce# => X"bc020000",
		16#37cf# => X"10000005",
		16#37d0# => X"85610030",
		16#37d1# => X"9c80ffff",
		16#37d2# => X"d4012030",
		16#37d3# => X"85610030",
		16#37d4# => X"9c210588",
		16#37d5# => X"8521fffc",
		16#37d6# => X"8441ffd4",
		16#37d7# => X"85c1ffd8",
		16#37d8# => X"8601ffdc",
		16#37d9# => X"8641ffe0",
		16#37da# => X"8681ffe4",
		16#37db# => X"86c1ffe8",
		16#37dc# => X"8701ffec",
		16#37dd# => X"8741fff0",
		16#37de# => X"8781fff4",
		16#37df# => X"44004800",
		16#37e0# => X"87c1fff8",
		16#37e1# => X"98e3000e",
		16#37e2# => X"bd870000",
		16#37e3# => X"13ffff1b",
		16#37e4# => X"9c80fffd",
		16#37e5# => X"9e010468",
		16#37e6# => X"e0422003",
		16#37e7# => X"85e30064",
		16#37e8# => X"85a3001c",
		16#37e9# => X"85830024",
		16#37ea# => X"9d610068",
		16#37eb# => X"9d000400",
		16#37ec# => X"dc011474",
		16#37ed# => X"84610028",
		16#37ee# => X"9c400000",
		16#37ef# => X"a8900000",
		16#37f0# => X"a8ae0000",
		16#37f1# => X"84c1002c",
		16#37f2# => X"d4017ccc",
		16#37f3# => X"dc013c76",
		16#37f4# => X"d4016c84",
		16#37f5# => X"d401648c",
		16#37f6# => X"d4015c68",
		16#37f7# => X"d4015c78",
		16#37f8# => X"d4014470",
		16#37f9# => X"d401447c",
		16#37fa# => X"07fffecc",
		16#37fb# => X"d4011480",
		16#37fc# => X"e58b1000",
		16#37fd# => X"10000008",
		16#37fe# => X"d4015830",
		16#37ff# => X"84610028",
		16#3800# => X"04001080",
		16#3801# => X"a8900000",
		16#3802# => X"e42b1000",
		16#3803# => X"100006fd",
		16#3804# => X"9c60ffff",
		16#3805# => X"94410474",
		16#3806# => X"a4420040",
		16#3807# => X"bc020000",
		16#3808# => X"13ffffcb",
		16#3809# => X"84810020",
		16#380a# => X"9444000c",
		16#380b# => X"a8420040",
		16#380c# => X"03ffffc7",
		16#380d# => X"dc04100c",
		16#380e# => X"04001180",
		16#380f# => X"84610028",
		16#3810# => X"03fffed4",
		16#3811# => X"84610020",
		16#3812# => X"85c1001c",
		16#3813# => X"03ffff2e",
		16#3814# => X"90ae0000",
		16#3815# => X"84610018",
		16#3816# => X"d401281c",
		16#3817# => X"a8630010",
		16#3818# => X"d801455b",
		16#3819# => X"d4011818",
		16#381a# => X"84810018",
		16#381b# => X"a4e40010",
		16#381c# => X"bc070000",
		16#381d# => X"0c000094",
		16#381e# => X"8441002c",
		16#381f# => X"84610018",
		16#3820# => X"a4e30040",
		16#3821# => X"bc070000",
		16#3822# => X"1000008f",
		16#3823# => X"8441002c",
		16#3824# => X"8481002c",
		16#3825# => X"99c40002",
		16#3826# => X"9c840004",
		16#3827# => X"d401202c",
		16#3828# => X"bd8e0000",
		16#3829# => X"1000043e",
		16#382a# => X"e0e07002",
		16#382b# => X"9d000001",
		16#382c# => X"e0e77004",
		16#382d# => X"b967005f",
		16#382e# => X"bd920000",
		16#382f# => X"10000005",
		16#3830# => X"84610018",
		16#3831# => X"9c80ff7f",
		16#3832# => X"e0632003",
		16#3833# => X"d4011818",
		16#3834# => X"e0e09002",
		16#3835# => X"e0e79004",
		16#3836# => X"bd870000",
		16#3837# => X"10000006",
		16#3838# => X"bc080001",
		16#3839# => X"bc0b0000",
		16#383a# => X"10000260",
		16#383b# => X"bc280000",
		16#383c# => X"bc080001",
		16#383d# => X"10000395",
		16#383e# => X"bc080002",
		16#383f# => X"10000384",
		16#3840# => X"9c410538",
		16#3841# => X"d4011040",
		16#3842# => X"a8620000",
		16#3843# => X"a44e0007",
		16#3844# => X"9c63ffff",
		16#3845# => X"9d020030",
		16#3846# => X"b9ce0043",
		16#3847# => X"bc2e0000",
		16#3848# => X"13fffffb",
		16#3849# => X"d8034000",
		16#384a# => X"d4011840",
		16#384b# => X"84610018",
		16#384c# => X"a4e30001",
		16#384d# => X"bc270000",
		16#384e# => X"10000410",
		16#384f# => X"bc280030",
		16#3850# => X"84810014",
		16#3851# => X"84410040",
		16#3852# => X"e3441002",
		16#3853# => X"e57a9000",
		16#3854# => X"10000003",
		16#3855# => X"d401d024",
		16#3856# => X"d4019024",
		16#3857# => X"9101055b",
		16#3858# => X"d4019044",
		16#3859# => X"bc080000",
		16#385a# => X"13ffff07",
		16#385b# => X"84410018",
		16#385c# => X"84810024",
		16#385d# => X"9c840001",
		16#385e# => X"03ffff02",
		16#385f# => X"d4012024",
		16#3860# => X"d801455b",
		16#3861# => X"d401281c",
		16#3862# => X"8441002c",
		16#3863# => X"8461002c",
		16#3864# => X"84420000",
		16#3865# => X"8481002c",
		16#3866# => X"d401104c",
		16#3867# => X"9c840008",
		16#3868# => X"84630004",
		16#3869# => X"8581004c",
		16#386a# => X"d4011850",
		16#386b# => X"a8ec0000",
		16#386c# => X"85610050",
		16#386d# => X"d401202c",
		16#386e# => X"a90b0000",
		16#386f# => X"e0670004",
		16#3870# => X"e0880004",
		16#3871# => X"04001da5",
		16#3872# => X"aa9e0000",
		16#3873# => X"bc2b0001",
		16#3874# => X"10000408",
		16#3875# => X"85a1004c",
		16#3876# => X"84a1004c",
		16#3877# => X"85610050",
		16#3878# => X"18400001",
		16#3879# => X"a8e50000",
		16#387a# => X"a90b0000",
		16#387b# => X"a84288d0",
		16#387c# => X"e0670004",
		16#387d# => X"e0880004",
		16#387e# => X"84a20000",
		16#387f# => X"84c20004",
		16#3880# => X"07fff717",
		16#3881# => X"15000000",
		16#3882# => X"bd8b0000",
		16#3883# => X"10000572",
		16#3884# => X"9c60002d",
		16#3885# => X"9101055b",
		16#3886# => X"18800001",
		16#3887# => X"bd5e0047",
		16#3888# => X"a884889a",
		16#3889# => X"10000005",
		16#388a# => X"d4012040",
		16#388b# => X"18400001",
		16#388c# => X"a8428896",
		16#388d# => X"d4011040",
		16#388e# => X"9c600003",
		16#388f# => X"84810018",
		16#3890# => X"9c40ff7f",
		16#3891# => X"d4011824",
		16#3892# => X"e0841003",
		16#3893# => X"ab430000",
		16#3894# => X"9c600000",
		16#3895# => X"d4012018",
		16#3896# => X"03ffffc3",
		16#3897# => X"d4011844",
		16#3898# => X"84810018",
		16#3899# => X"a8840008",
		16#389a# => X"03fffeb2",
		16#389b# => X"d4012018",
		16#389c# => X"8441002c",
		16#389d# => X"d401281c",
		16#389e# => X"84a20000",
		16#389f# => X"9c420004",
		16#38a0# => X"9c600001",
		16#38a1# => X"9c800000",
		16#38a2# => X"d401102c",
		16#38a3# => X"9c410510",
		16#38a4# => X"d4011824",
		16#38a5# => X"d8012d10",
		16#38a6# => X"d801255b",
		16#38a7# => X"ab430000",
		16#38a8# => X"03fffeb6",
		16#38a9# => X"d4011040",
		16#38aa# => X"84810018",
		16#38ab# => X"d401281c",
		16#38ac# => X"a4e40010",
		16#38ad# => X"bc070000",
		16#38ae# => X"13ffff71",
		16#38af# => X"d801455b",
		16#38b0# => X"8441002c",
		16#38b1# => X"85c20000",
		16#38b2# => X"9c420004",
		16#38b3# => X"03ffff75",
		16#38b4# => X"d401102c",
		16#38b5# => X"bc280000",
		16#38b6# => X"13fffe96",
		16#38b7# => X"15000000",
		16#38b8# => X"03fffe94",
		16#38b9# => X"9d000020",
		16#38ba# => X"84810018",
		16#38bb# => X"a8840001",
		16#38bc# => X"03fffe90",
		16#38bd# => X"d4012018",
		16#38be# => X"03fffe8e",
		16#38bf# => X"9d00002b",
		16#38c0# => X"84610018",
		16#38c1# => X"a8630080",
		16#38c2# => X"03fffe8a",
		16#38c3# => X"d4011818",
		16#38c4# => X"9c400000",
		16#38c5# => X"9c9effd0",
		16#38c6# => X"b8620003",
		16#38c7# => X"e0421000",
		16#38c8# => X"93c50000",
		16#38c9# => X"e0421800",
		16#38ca# => X"e0441000",
		16#38cb# => X"9c9effd0",
		16#38cc# => X"bca40009",
		16#38cd# => X"13fffff9",
		16#38ce# => X"9ca50001",
		16#38cf# => X"03fffe7f",
		16#38d0# => X"d4011034",
		16#38d1# => X"93c50000",
		16#38d2# => X"bc1e002a",
		16#38d3# => X"1000061d",
		16#38d4# => X"9ca50001",
		16#38d5# => X"9c9effd0",
		16#38d6# => X"bca40009",
		16#38d7# => X"0c00000b",
		16#38d8# => X"9e400000",
		16#38d9# => X"b8520003",
		16#38da# => X"e2529000",
		16#38db# => X"93c50000",
		16#38dc# => X"e2521000",
		16#38dd# => X"e2522000",
		16#38de# => X"9c9effd0",
		16#38df# => X"bca40009",
		16#38e0# => X"13fffff9",
		16#38e1# => X"9ca50001",
		16#38e2# => X"bd720000",
		16#38e3# => X"13fffe6c",
		16#38e4# => X"9c7effe0",
		16#38e5# => X"03fffe6a",
		16#38e6# => X"9e40ffff",
		16#38e7# => X"84410018",
		16#38e8# => X"a8420040",
		16#38e9# => X"03fffe63",
		16#38ea# => X"d4011018",
		16#38eb# => X"84610018",
		16#38ec# => X"a8630010",
		16#38ed# => X"03fffe5f",
		16#38ee# => X"d4011818",
		16#38ef# => X"84410018",
		16#38f0# => X"d401281c",
		16#38f1# => X"a4a20010",
		16#38f2# => X"bc050000",
		16#38f3# => X"10000451",
		16#38f4# => X"d801455b",
		16#38f5# => X"8461002c",
		16#38f6# => X"84810030",
		16#38f7# => X"84430000",
		16#38f8# => X"9c630004",
		16#38f9# => X"d401182c",
		16#38fa# => X"03fffe1e",
		16#38fb# => X"d4022000",
		16#38fc# => X"8481002c",
		16#38fd# => X"84410018",
		16#38fe# => X"85c40000",
		16#38ff# => X"a8420002",
		16#3900# => X"9c600030",
		16#3901# => X"e0e07002",
		16#3902# => X"d4011018",
		16#3903# => X"d8011d58",
		16#3904# => X"8441002c",
		16#3905# => X"18600001",
		16#3906# => X"e0e77004",
		16#3907# => X"9c800078",
		16#3908# => X"9c420004",
		16#3909# => X"a86388b7",
		16#390a# => X"b967005f",
		16#390b# => X"d401281c",
		16#390c# => X"d8012559",
		16#390d# => X"d401102c",
		16#390e# => X"d401185c",
		16#390f# => X"9d000002",
		16#3910# => X"9fc00078",
		16#3911# => X"9c400000",
		16#3912# => X"03ffff1c",
		16#3913# => X"d801155b",
		16#3914# => X"9c800000",
		16#3915# => X"8441002c",
		16#3916# => X"d801255b",
		16#3917# => X"d401281c",
		16#3918# => X"84620000",
		16#3919# => X"9dc20004",
		16#391a# => X"bc230000",
		16#391b# => X"0c00053b",
		16#391c# => X"d4011840",
		16#391d# => X"bd920000",
		16#391e# => X"10000518",
		16#391f# => X"84610040",
		16#3920# => X"9c800000",
		16#3921# => X"040014ea",
		16#3922# => X"a8b20000",
		16#3923# => X"bc2b0000",
		16#3924# => X"0c000597",
		16#3925# => X"84410040",
		16#3926# => X"e34b1002",
		16#3927# => X"e5ba9000",
		16#3928# => X"100004ad",
		16#3929# => X"ac5affff",
		16#392a# => X"9c600000",
		16#392b# => X"d4019024",
		16#392c# => X"9101055b",
		16#392d# => X"ab520000",
		16#392e# => X"d401702c",
		16#392f# => X"03ffff2a",
		16#3930# => X"d4011844",
		16#3931# => X"18600001",
		16#3932# => X"84810018",
		16#3933# => X"a86388b7",
		16#3934# => X"a4e40010",
		16#3935# => X"d401281c",
		16#3936# => X"d801455b",
		16#3937# => X"bc070000",
		16#3938# => X"0c00003c",
		16#3939# => X"d401185c",
		16#393a# => X"84610018",
		16#393b# => X"a4e30040",
		16#393c# => X"bc070000",
		16#393d# => X"10000038",
		16#393e# => X"8441002c",
		16#393f# => X"8481002c",
		16#3940# => X"85c40000",
		16#3941# => X"9c840004",
		16#3942# => X"a5ceffff",
		16#3943# => X"e0e07002",
		16#3944# => X"e0e77004",
		16#3945# => X"b967005f",
		16#3946# => X"bc0b0000",
		16#3947# => X"10000036",
		16#3948# => X"d401202c",
		16#3949# => X"84610018",
		16#394a# => X"a5030001",
		16#394b# => X"bc080000",
		16#394c# => X"10000031",
		16#394d# => X"9c800030",
		16#394e# => X"a8630002",
		16#394f# => X"d8012558",
		16#3950# => X"d801f559",
		16#3951# => X"d4011818",
		16#3952# => X"9d600001",
		16#3953# => X"03ffffbe",
		16#3954# => X"9d000002",
		16#3955# => X"84810018",
		16#3956# => X"a8840010",
		16#3957# => X"03fffdf5",
		16#3958# => X"d4012018",
		16#3959# => X"84610018",
		16#395a# => X"d401281c",
		16#395b# => X"a8630010",
		16#395c# => X"d4011818",
		16#395d# => X"84810018",
		16#395e# => X"a4e40010",
		16#395f# => X"bc070000",
		16#3960# => X"100002b7",
		16#3961# => X"84610018",
		16#3962# => X"8441002c",
		16#3963# => X"9d000001",
		16#3964# => X"85c20000",
		16#3965# => X"9c420004",
		16#3966# => X"e0e07002",
		16#3967# => X"d401102c",
		16#3968# => X"e0e77004",
		16#3969# => X"03ffffa8",
		16#396a# => X"b967005f",
		16#396b# => X"18600001",
		16#396c# => X"84810018",
		16#396d# => X"a86388a6",
		16#396e# => X"a4e40010",
		16#396f# => X"d401281c",
		16#3970# => X"d801455b",
		16#3971# => X"bc070000",
		16#3972# => X"13ffffc8",
		16#3973# => X"d401185c",
		16#3974# => X"8441002c",
		16#3975# => X"85c20000",
		16#3976# => X"9c420004",
		16#3977# => X"e0e07002",
		16#3978# => X"e0e77004",
		16#3979# => X"b967005f",
		16#397a# => X"bc0b0000",
		16#397b# => X"0fffffce",
		16#397c# => X"d401102c",
		16#397d# => X"03ffff94",
		16#397e# => X"9d000002",
		16#397f# => X"84810018",
		16#3980# => X"d401281c",
		16#3981# => X"a8840010",
		16#3982# => X"d4012018",
		16#3983# => X"84410018",
		16#3984# => X"a5020010",
		16#3985# => X"bc080000",
		16#3986# => X"1000029e",
		16#3987# => X"84810018",
		16#3988# => X"8461002c",
		16#3989# => X"9d000000",
		16#398a# => X"85c30000",
		16#398b# => X"9c630004",
		16#398c# => X"e0e07002",
		16#398d# => X"d401182c",
		16#398e# => X"e0e77004",
		16#398f# => X"03ffff82",
		16#3990# => X"b967005f",
		16#3991# => X"03fffff2",
		16#3992# => X"d401281c",
		16#3993# => X"03ffffca",
		16#3994# => X"d401281c",
		16#3995# => X"9f160008",
		16#3996# => X"86410540",
		16#3997# => X"8601053c",
		16#3998# => X"9041055b",
		16#3999# => X"bc020000",
		16#399a# => X"1000000f",
		16#399b# => X"bc1c0000",
		16#399c# => X"9e100001",
		16#399d# => X"9e520001",
		16#399e# => X"9c81055b",
		16#399f# => X"9c400001",
		16#39a0# => X"d4162000",
		16#39a1# => X"d4161004",
		16#39a2# => X"d4019540",
		16#39a3# => X"bd500007",
		16#39a4# => X"100001d0",
		16#39a5# => X"d401853c",
		16#39a6# => X"aad80000",
		16#39a7# => X"9f180008",
		16#39a8# => X"bc1c0000",
		16#39a9# => X"1000000f",
		16#39aa# => X"8441003c",
		16#39ab# => X"9e100001",
		16#39ac# => X"9e520002",
		16#39ad# => X"9c610558",
		16#39ae# => X"9c800002",
		16#39af# => X"d4161800",
		16#39b0# => X"d4162004",
		16#39b1# => X"d4019540",
		16#39b2# => X"bd500007",
		16#39b3# => X"100001cc",
		16#39b4# => X"d401853c",
		16#39b5# => X"aad80000",
		16#39b6# => X"9f180008",
		16#39b7# => X"8441003c",
		16#39b8# => X"bc220080",
		16#39b9# => X"0c0000ee",
		16#39ba# => X"84610034",
		16#39bb# => X"84610044",
		16#39bc# => X"e043d002",
		16#39bd# => X"bda20000",
		16#39be# => X"1000002e",
		16#39bf# => X"bda20010",
		16#39c0# => X"100003c5",
		16#39c1# => X"15000000",
		16#39c2# => X"1a800001",
		16#39c3# => X"9dc00010",
		16#39c4# => X"aa948a3c",
		16#39c5# => X"87010028",
		16#39c6# => X"00000007",
		16#39c7# => X"87810020",
		16#39c8# => X"9ed60008",
		16#39c9# => X"9c42fff0",
		16#39ca# => X"bd420010",
		16#39cb# => X"0c000017",
		16#39cc# => X"9cb60008",
		16#39cd# => X"9e100001",
		16#39ce# => X"9e520010",
		16#39cf# => X"d416a000",
		16#39d0# => X"d4167004",
		16#39d1# => X"d4019540",
		16#39d2# => X"bd500007",
		16#39d3# => X"0ffffff5",
		16#39d4# => X"d401853c",
		16#39d5# => X"a8780000",
		16#39d6# => X"a89c0000",
		16#39d7# => X"04001d3f",
		16#39d8# => X"9ca10538",
		16#39d9# => X"bc2b0000",
		16#39da# => X"13fffdf1",
		16#39db# => X"9c42fff0",
		16#39dc# => X"9ca104d8",
		16#39dd# => X"9ec104d0",
		16#39de# => X"86410540",
		16#39df# => X"bd420010",
		16#39e0# => X"13ffffed",
		16#39e1# => X"8601053c",
		16#39e2# => X"9e100001",
		16#39e3# => X"e2521000",
		16#39e4# => X"d416a000",
		16#39e5# => X"d4161004",
		16#39e6# => X"d4019540",
		16#39e7# => X"bd500007",
		16#39e8# => X"10000181",
		16#39e9# => X"d401853c",
		16#39ea# => X"9f050008",
		16#39eb# => X"aac50000",
		16#39ec# => X"84810018",
		16#39ed# => X"a4440100",
		16#39ee# => X"bc220000",
		16#39ef# => X"10000054",
		16#39f0# => X"bdbe0065",
		16#39f1# => X"9e100001",
		16#39f2# => X"e252d000",
		16#39f3# => X"84410040",
		16#39f4# => X"d416d004",
		16#39f5# => X"d4161000",
		16#39f6# => X"d4019540",
		16#39f7# => X"bdb00007",
		16#39f8# => X"0c00010c",
		16#39f9# => X"d401853c",
		16#39fa# => X"84810018",
		16#39fb# => X"a4440004",
		16#39fc# => X"bc220000",
		16#39fd# => X"0c000039",
		16#39fe# => X"84410024",
		16#39ff# => X"84410034",
		16#3a00# => X"84610024",
		16#3a01# => X"e1c21802",
		16#3a02# => X"bd4e0000",
		16#3a03# => X"0c000032",
		16#3a04# => X"bdae0010",
		16#3a05# => X"10000468",
		16#3a06# => X"15000000",
		16#3a07# => X"1a800001",
		16#3a08# => X"8601053c",
		16#3a09# => X"aa948a4c",
		16#3a0a# => X"9ec00010",
		16#3a0b# => X"84410028",
		16#3a0c# => X"00000006",
		16#3a0d# => X"87410020",
		16#3a0e# => X"9dcefff0",
		16#3a0f# => X"bd4e0010",
		16#3a10# => X"0c000016",
		16#3a11# => X"9f180008",
		16#3a12# => X"9e100001",
		16#3a13# => X"9e520010",
		16#3a14# => X"d418a000",
		16#3a15# => X"d418b004",
		16#3a16# => X"d4019540",
		16#3a17# => X"bd500007",
		16#3a18# => X"0ffffff6",
		16#3a19# => X"d401853c",
		16#3a1a# => X"a8620000",
		16#3a1b# => X"a89a0000",
		16#3a1c# => X"04001cfa",
		16#3a1d# => X"9ca10538",
		16#3a1e# => X"bc2b0000",
		16#3a1f# => X"13fffdac",
		16#3a20# => X"9dcefff0",
		16#3a21# => X"9f0104d0",
		16#3a22# => X"86410540",
		16#3a23# => X"bd4e0010",
		16#3a24# => X"13ffffee",
		16#3a25# => X"8601053c",
		16#3a26# => X"9e100001",
		16#3a27# => X"e24e9000",
		16#3a28# => X"d418a000",
		16#3a29# => X"d4187004",
		16#3a2a# => X"d4019540",
		16#3a2b# => X"bdb00007",
		16#3a2c# => X"10000009",
		16#3a2d# => X"d401853c",
		16#3a2e# => X"84610028",
		16#3a2f# => X"84810020",
		16#3a30# => X"04001ce6",
		16#3a31# => X"9ca10538",
		16#3a32# => X"bc2b0000",
		16#3a33# => X"13fffd98",
		16#3a34# => X"86410540",
		16#3a35# => X"84410024",
		16#3a36# => X"84810034",
		16#3a37# => X"e5622000",
		16#3a38# => X"10000003",
		16#3a39# => X"84610030",
		16#3a3a# => X"a8440000",
		16#3a3b# => X"bc120000",
		16#3a3c# => X"e0631000",
		16#3a3d# => X"0c00009c",
		16#3a3e# => X"d4011830",
		16#3a3f# => X"9c800000",
		16#3a40# => X"9ec104d0",
		16#3a41# => X"03fffcd7",
		16#3a42# => X"d401253c",
		16#3a43# => X"100000ca",
		16#3a44# => X"84410038",
		16#3a45# => X"84a1004c",
		16#3a46# => X"85810050",
		16#3a47# => X"18600001",
		16#3a48# => X"a8e50000",
		16#3a49# => X"a86388d0",
		16#3a4a# => X"a90c0000",
		16#3a4b# => X"84a30000",
		16#3a4c# => X"84c30004",
		16#3a4d# => X"e0670004",
		16#3a4e# => X"e0880004",
		16#3a4f# => X"07fff4d0",
		16#3a50# => X"15000000",
		16#3a51# => X"bc0b0000",
		16#3a52# => X"0c000138",
		16#3a53# => X"85c10554",
		16#3a54# => X"18a00001",
		16#3a55# => X"9e100001",
		16#3a56# => X"9e520001",
		16#3a57# => X"a8a5842b",
		16#3a58# => X"9c800001",
		16#3a59# => X"d4162800",
		16#3a5a# => X"d4162004",
		16#3a5b# => X"d4019540",
		16#3a5c# => X"bdb00007",
		16#3a5d# => X"0c00032c",
		16#3a5e# => X"d401853c",
		16#3a5f# => X"84a10554",
		16#3a60# => X"84410038",
		16#3a61# => X"e5851000",
		16#3a62# => X"10000006",
		16#3a63# => X"84610018",
		16#3a64# => X"a4a30001",
		16#3a65# => X"bc050000",
		16#3a66# => X"13ffff95",
		16#3a67# => X"84810018",
		16#3a68# => X"8601053c",
		16#3a69# => X"84810054",
		16#3a6a# => X"9e100001",
		16#3a6b# => X"e2522000",
		16#3a6c# => X"84410048",
		16#3a6d# => X"d4182004",
		16#3a6e# => X"d4181000",
		16#3a6f# => X"d4019540",
		16#3a70# => X"bd500007",
		16#3a71# => X"100003ac",
		16#3a72# => X"d401853c",
		16#3a73# => X"9cb80008",
		16#3a74# => X"84610038",
		16#3a75# => X"9dc3ffff",
		16#3a76# => X"bdae0000",
		16#3a77# => X"100003af",
		16#3a78# => X"bd4e0010",
		16#3a79# => X"0c0001f6",
		16#3a7a# => X"1a800001",
		16#3a7b# => X"8601053c",
		16#3a7c# => X"aa948a3c",
		16#3a7d# => X"9ec00010",
		16#3a7e# => X"84410028",
		16#3a7f# => X"00000008",
		16#3a80# => X"87410020",
		16#3a81# => X"9ca50008",
		16#3a82# => X"9f050008",
		16#3a83# => X"9dcefff0",
		16#3a84# => X"bd4e0010",
		16#3a85# => X"0c0001ed",
		16#3a86# => X"15000000",
		16#3a87# => X"9e100001",
		16#3a88# => X"9e520010",
		16#3a89# => X"d405a000",
		16#3a8a# => X"d405b004",
		16#3a8b# => X"d4019540",
		16#3a8c# => X"bd500007",
		16#3a8d# => X"0ffffff4",
		16#3a8e# => X"d401853c",
		16#3a8f# => X"a8620000",
		16#3a90# => X"a89a0000",
		16#3a91# => X"04001c85",
		16#3a92# => X"9ca10538",
		16#3a93# => X"bc2b0000",
		16#3a94# => X"13fffd37",
		16#3a95# => X"9f0104d8",
		16#3a96# => X"9ca104d0",
		16#3a97# => X"86410540",
		16#3a98# => X"03ffffeb",
		16#3a99# => X"8601053c",
		16#3a9a# => X"100000cc",
		16#3a9b# => X"9c410538",
		16#3a9c# => X"84410018",
		16#3a9d# => X"a4e20001",
		16#3a9e# => X"bc070000",
		16#3a9f# => X"10000121",
		16#3aa0# => X"9c610538",
		16#3aa1# => X"9c600030",
		16#3aa2# => X"9c810537",
		16#3aa3# => X"d8011d37",
		16#3aa4# => X"87410064",
		16#3aa5# => X"03fffdae",
		16#3aa6# => X"d4012040",
		16#3aa7# => X"84810024",
		16#3aa8# => X"e1c32002",
		16#3aa9# => X"bd4e0000",
		16#3aaa# => X"0c000186",
		16#3aab# => X"bdae0010",
		16#3aac# => X"1000040b",
		16#3aad# => X"15000000",
		16#3aae# => X"1a800001",
		16#3aaf# => X"9f000010",
		16#3ab0# => X"aa948a3c",
		16#3ab1# => X"84410028",
		16#3ab2# => X"00000007",
		16#3ab3# => X"87810020",
		16#3ab4# => X"9ed60008",
		16#3ab5# => X"9dcefff0",
		16#3ab6# => X"bd4e0010",
		16#3ab7# => X"0c000017",
		16#3ab8# => X"9d160008",
		16#3ab9# => X"9e100001",
		16#3aba# => X"9e520010",
		16#3abb# => X"d416a000",
		16#3abc# => X"d416c004",
		16#3abd# => X"d4019540",
		16#3abe# => X"bd500007",
		16#3abf# => X"0ffffff5",
		16#3ac0# => X"d401853c",
		16#3ac1# => X"a8620000",
		16#3ac2# => X"a89c0000",
		16#3ac3# => X"04001c53",
		16#3ac4# => X"9ca10538",
		16#3ac5# => X"bc2b0000",
		16#3ac6# => X"13fffd05",
		16#3ac7# => X"9dcefff0",
		16#3ac8# => X"9d0104d8",
		16#3ac9# => X"9ec104d0",
		16#3aca# => X"86410540",
		16#3acb# => X"bd4e0010",
		16#3acc# => X"13ffffed",
		16#3acd# => X"8601053c",
		16#3ace# => X"9e100001",
		16#3acf# => X"e2527000",
		16#3ad0# => X"d416a000",
		16#3ad1# => X"d4167004",
		16#3ad2# => X"d4019540",
		16#3ad3# => X"bd500007",
		16#3ad4# => X"1000017f",
		16#3ad5# => X"d401853c",
		16#3ad6# => X"9f080008",
		16#3ad7# => X"03fffee4",
		16#3ad8# => X"aac80000",
		16#3ad9# => X"84610028",
		16#3ada# => X"84810020",
		16#3adb# => X"04001c3b",
		16#3adc# => X"9ca10538",
		16#3add# => X"bc2b0000",
		16#3ade# => X"0fffff62",
		16#3adf# => X"9c800000",
		16#3ae0# => X"03fffcec",
		16#3ae1# => X"84610020",
		16#3ae2# => X"9e100001",
		16#3ae3# => X"84410040",
		16#3ae4# => X"d4161000",
		16#3ae5# => X"d4167004",
		16#3ae6# => X"d4015d40",
		16#3ae7# => X"d401853c",
		16#3ae8# => X"bdb00007",
		16#3ae9# => X"0c000388",
		16#3aea# => X"a84e0000",
		16#3aeb# => X"84610054",
		16#3aec# => X"9e100001",
		16#3aed# => X"e16b1800",
		16#3aee# => X"84810048",
		16#3aef# => X"d4181804",
		16#3af0# => X"d4182000",
		16#3af1# => X"d4015d40",
		16#3af2# => X"bd500007",
		16#3af3# => X"10000391",
		16#3af4# => X"d401853c",
		16#3af5# => X"9f180008",
		16#3af6# => X"84610038",
		16#3af7# => X"86410540",
		16#3af8# => X"e1c37002",
		16#3af9# => X"8601053c",
		16#3afa# => X"84810040",
		16#3afb# => X"9e100001",
		16#3afc# => X"e1041000",
		16#3afd# => X"e2527000",
		16#3afe# => X"d4184000",
		16#3aff# => X"d4187004",
		16#3b00# => X"d4019540",
		16#3b01# => X"bd500007",
		16#3b02# => X"0c000281",
		16#3b03# => X"d401853c",
		16#3b04# => X"84610028",
		16#3b05# => X"84810020",
		16#3b06# => X"04001c10",
		16#3b07# => X"9ca10538",
		16#3b08# => X"bc2b0000",
		16#3b09# => X"13fffcc2",
		16#3b0a# => X"9f0104d0",
		16#3b0b# => X"03fffeef",
		16#3b0c# => X"86410540",
		16#3b0d# => X"bd420001",
		16#3b0e# => X"0c000040",
		16#3b0f# => X"84610018",
		16#3b10# => X"9e100001",
		16#3b11# => X"9e520001",
		16#3b12# => X"84810040",
		16#3b13# => X"9c400001",
		16#3b14# => X"d4162000",
		16#3b15# => X"d4161004",
		16#3b16# => X"d4019540",
		16#3b17# => X"bd500007",
		16#3b18# => X"1000011a",
		16#3b19# => X"d401853c",
		16#3b1a# => X"9dd80008",
		16#3b1b# => X"84610054",
		16#3b1c# => X"9e100001",
		16#3b1d# => X"e2521800",
		16#3b1e# => X"84810048",
		16#3b1f# => X"d4181804",
		16#3b20# => X"d4182000",
		16#3b21# => X"d4019540",
		16#3b22# => X"bd500007",
		16#3b23# => X"1000011a",
		16#3b24# => X"d401853c",
		16#3b25# => X"9f4e0008",
		16#3b26# => X"84a1004c",
		16#3b27# => X"85810050",
		16#3b28# => X"18400001",
		16#3b29# => X"a8e50000",
		16#3b2a# => X"a90c0000",
		16#3b2b# => X"a84288d0",
		16#3b2c# => X"e0670004",
		16#3b2d# => X"e0880004",
		16#3b2e# => X"84a20000",
		16#3b2f# => X"84c20004",
		16#3b30# => X"07fff40d",
		16#3b31# => X"15000000",
		16#3b32# => X"bc2b0000",
		16#3b33# => X"0c0000c0",
		16#3b34# => X"84410038",
		16#3b35# => X"84610038",
		16#3b36# => X"84810040",
		16#3b37# => X"9d03ffff",
		16#3b38# => X"9e100001",
		16#3b39# => X"9ca40001",
		16#3b3a# => X"e2524000",
		16#3b3b# => X"d40e2800",
		16#3b3c# => X"d40e4004",
		16#3b3d# => X"d4019540",
		16#3b3e# => X"bd500007",
		16#3b3f# => X"1000001c",
		16#3b40# => X"d401853c",
		16#3b41# => X"9f1a0008",
		16#3b42# => X"84410058",
		16#3b43# => X"9e100001",
		16#3b44# => X"e2521000",
		16#3b45# => X"9c610544",
		16#3b46# => X"d41a1004",
		16#3b47# => X"d41a1800",
		16#3b48# => X"d4019540",
		16#3b49# => X"bdb00007",
		16#3b4a# => X"13fffeb0",
		16#3b4b# => X"d401853c",
		16#3b4c# => X"03ffffb9",
		16#3b4d# => X"84610028",
		16#3b4e# => X"a4a30001",
		16#3b4f# => X"bc050000",
		16#3b50# => X"0fffffc0",
		16#3b51# => X"84610040",
		16#3b52# => X"9e100001",
		16#3b53# => X"9e520001",
		16#3b54# => X"9c800001",
		16#3b55# => X"d4161800",
		16#3b56# => X"d4162004",
		16#3b57# => X"d4019540",
		16#3b58# => X"bd500007",
		16#3b59# => X"0c00029f",
		16#3b5a# => X"d401853c",
		16#3b5b# => X"84610028",
		16#3b5c# => X"84810020",
		16#3b5d# => X"04001bb9",
		16#3b5e# => X"9ca10538",
		16#3b5f# => X"bc2b0000",
		16#3b60# => X"13fffc6b",
		16#3b61# => X"9f0104d8",
		16#3b62# => X"9f4104d0",
		16#3b63# => X"86410540",
		16#3b64# => X"03ffffde",
		16#3b65# => X"8601053c",
		16#3b66# => X"ab4b0000",
		16#3b67# => X"03fffcec",
		16#3b68# => X"d4011040",
		16#3b69# => X"84610028",
		16#3b6a# => X"84810020",
		16#3b6b# => X"04001bab",
		16#3b6c# => X"9ca10538",
		16#3b6d# => X"bc2b0000",
		16#3b6e# => X"13fffc5d",
		16#3b6f# => X"9f0104d8",
		16#3b70# => X"9ec104d0",
		16#3b71# => X"86410540",
		16#3b72# => X"03fffe7a",
		16#3b73# => X"8601053c",
		16#3b74# => X"84610028",
		16#3b75# => X"84810020",
		16#3b76# => X"04001ba0",
		16#3b77# => X"9ca10538",
		16#3b78# => X"bc2b0000",
		16#3b79# => X"13fffc52",
		16#3b7a# => X"9f0104d8",
		16#3b7b# => X"9ec104d0",
		16#3b7c# => X"86410540",
		16#3b7d# => X"03fffe2b",
		16#3b7e# => X"8601053c",
		16#3b7f# => X"84610028",
		16#3b80# => X"84810020",
		16#3b81# => X"04001b95",
		16#3b82# => X"9ca10538",
		16#3b83# => X"bc2b0000",
		16#3b84# => X"13fffc47",
		16#3b85# => X"9f0104d8",
		16#3b86# => X"9ec104d0",
		16#3b87# => X"86410540",
		16#3b88# => X"03fffe2f",
		16#3b89# => X"8601053c",
		16#3b8a# => X"bd4e0000",
		16#3b8b# => X"0c000207",
		16#3b8c# => X"84410038",
		16#3b8d# => X"e58e1000",
		16#3b8e# => X"13ffff54",
		16#3b8f# => X"e16e9000",
		16#3b90# => X"9e100001",
		16#3b91# => X"e2521000",
		16#3b92# => X"84610040",
		16#3b93# => X"d4161004",
		16#3b94# => X"d4161800",
		16#3b95# => X"d4019540",
		16#3b96# => X"bdb00007",
		16#3b97# => X"0c0002f6",
		16#3b98# => X"d401853c",
		16#3b99# => X"84810038",
		16#3b9a# => X"e1ce2002",
		16#3b9b# => X"bdae0000",
		16#3b9c# => X"100001d7",
		16#3b9d# => X"bd4e0010",
		16#3b9e# => X"0c0001c1",
		16#3b9f# => X"1a800001",
		16#3ba0# => X"a8b80000",
		16#3ba1# => X"8601053c",
		16#3ba2# => X"aa948a3c",
		16#3ba3# => X"9ec00010",
		16#3ba4# => X"84410028",
		16#3ba5# => X"00000008",
		16#3ba6# => X"87410020",
		16#3ba7# => X"9ca50008",
		16#3ba8# => X"9f050008",
		16#3ba9# => X"9dcefff0",
		16#3baa# => X"bd4e0010",
		16#3bab# => X"0c0001b8",
		16#3bac# => X"15000000",
		16#3bad# => X"9e100001",
		16#3bae# => X"9e520010",
		16#3baf# => X"d405a000",
		16#3bb0# => X"d405b004",
		16#3bb1# => X"d4019540",
		16#3bb2# => X"bd500007",
		16#3bb3# => X"0ffffff4",
		16#3bb4# => X"d401853c",
		16#3bb5# => X"a8620000",
		16#3bb6# => X"a89a0000",
		16#3bb7# => X"04001b5f",
		16#3bb8# => X"9ca10538",
		16#3bb9# => X"bc2b0000",
		16#3bba# => X"13fffc11",
		16#3bbb# => X"9f0104d8",
		16#3bbc# => X"9ca104d0",
		16#3bbd# => X"86410540",
		16#3bbe# => X"03ffffeb",
		16#3bbf# => X"8601053c",
		16#3bc0# => X"ab480000",
		16#3bc1# => X"03fffc92",
		16#3bc2# => X"d4011840",
		16#3bc3# => X"9c610538",
		16#3bc4# => X"8481005c",
		16#3bc5# => X"d4011840",
		16#3bc6# => X"a44e000f",
		16#3bc7# => X"9c63ffff",
		16#3bc8# => X"e0441000",
		16#3bc9# => X"b9ce0044",
		16#3bca# => X"8c420000",
		16#3bcb# => X"bc2e0000",
		16#3bcc# => X"13fffffa",
		16#3bcd# => X"d8031000",
		16#3bce# => X"84810014",
		16#3bcf# => X"d4011840",
		16#3bd0# => X"03fffc83",
		16#3bd1# => X"e3441802",
		16#3bd2# => X"bc4e0009",
		16#3bd3# => X"0c00000e",
		16#3bd4# => X"9e010538",
		16#3bd5# => X"a86e0000",
		16#3bd6# => X"9c80000a",
		16#3bd7# => X"04002399",
		16#3bd8# => X"9e10ffff",
		16#3bd9# => X"9d6b0030",
		16#3bda# => X"a86e0000",
		16#3bdb# => X"9c80000a",
		16#3bdc# => X"07ffe9f0",
		16#3bdd# => X"d8105800",
		16#3bde# => X"bc4b0009",
		16#3bdf# => X"13fffff6",
		16#3be0# => X"a9cb0000",
		16#3be1# => X"9e10ffff",
		16#3be2# => X"84410014",
		16#3be3# => X"9dce0030",
		16#3be4# => X"d4018040",
		16#3be5# => X"e3428002",
		16#3be6# => X"03fffc6d",
		16#3be7# => X"d8107000",
		16#3be8# => X"84610028",
		16#3be9# => X"84810020",
		16#3bea# => X"04001b2c",
		16#3beb# => X"9ca10538",
		16#3bec# => X"bc2b0000",
		16#3bed# => X"13fffbde",
		16#3bee# => X"9f0104d8",
		16#3bef# => X"9ec104d0",
		16#3bf0# => X"86410540",
		16#3bf1# => X"03fffda7",
		16#3bf2# => X"8601053c",
		16#3bf3# => X"9ec2ffff",
		16#3bf4# => X"bd560000",
		16#3bf5# => X"0c000225",
		16#3bf6# => X"bdb60010",
		16#3bf7# => X"10000051",
		16#3bf8# => X"1a800001",
		16#3bf9# => X"9f000010",
		16#3bfa# => X"aa948a3c",
		16#3bfb# => X"84410028",
		16#3bfc# => X"00000008",
		16#3bfd# => X"87810020",
		16#3bfe# => X"9dce0008",
		16#3bff# => X"9f4e0008",
		16#3c00# => X"9ed6fff0",
		16#3c01# => X"bd560010",
		16#3c02# => X"0c000047",
		16#3c03# => X"15000000",
		16#3c04# => X"9e100001",
		16#3c05# => X"9e520010",
		16#3c06# => X"d40ea000",
		16#3c07# => X"d40ec004",
		16#3c08# => X"d4019540",
		16#3c09# => X"bd500007",
		16#3c0a# => X"0ffffff4",
		16#3c0b# => X"d401853c",
		16#3c0c# => X"a8620000",
		16#3c0d# => X"a89c0000",
		16#3c0e# => X"04001b08",
		16#3c0f# => X"9ca10538",
		16#3c10# => X"bc2b0000",
		16#3c11# => X"13fffbba",
		16#3c12# => X"9f4104d8",
		16#3c13# => X"9dc104d0",
		16#3c14# => X"86410540",
		16#3c15# => X"03ffffeb",
		16#3c16# => X"8601053c",
		16#3c17# => X"a4e30040",
		16#3c18# => X"bc070000",
		16#3c19# => X"10000136",
		16#3c1a# => X"8441002c",
		16#3c1b# => X"8481002c",
		16#3c1c# => X"9d000001",
		16#3c1d# => X"85c40000",
		16#3c1e# => X"9c840004",
		16#3c1f# => X"a5ceffff",
		16#3c20# => X"d401202c",
		16#3c21# => X"e0e07002",
		16#3c22# => X"03fffcef",
		16#3c23# => X"b967005f",
		16#3c24# => X"a5640040",
		16#3c25# => X"bc0b0000",
		16#3c26# => X"10000131",
		16#3c27# => X"8461002c",
		16#3c28# => X"8441002c",
		16#3c29# => X"85c20000",
		16#3c2a# => X"9c420004",
		16#3c2b# => X"a5ceffff",
		16#3c2c# => X"d401102c",
		16#3c2d# => X"e0e07002",
		16#3c2e# => X"03fffce3",
		16#3c2f# => X"b967005f",
		16#3c30# => X"03fffd8b",
		16#3c31# => X"9f160008",
		16#3c32# => X"84610028",
		16#3c33# => X"84810020",
		16#3c34# => X"04001ae2",
		16#3c35# => X"9ca10538",
		16#3c36# => X"bc2b0000",
		16#3c37# => X"13fffb94",
		16#3c38# => X"9dc104d8",
		16#3c39# => X"9f0104d0",
		16#3c3a# => X"86410540",
		16#3c3b# => X"03fffee0",
		16#3c3c# => X"8601053c",
		16#3c3d# => X"84610028",
		16#3c3e# => X"84810020",
		16#3c3f# => X"04001ad7",
		16#3c40# => X"9ca10538",
		16#3c41# => X"bc2b0000",
		16#3c42# => X"13fffb89",
		16#3c43# => X"9f4104d8",
		16#3c44# => X"9dc104d0",
		16#3c45# => X"86410540",
		16#3c46# => X"03fffee0",
		16#3c47# => X"8601053c",
		16#3c48# => X"aa948a3c",
		16#3c49# => X"9e100001",
		16#3c4a# => X"e252b000",
		16#3c4b# => X"d40ea000",
		16#3c4c# => X"d40eb004",
		16#3c4d# => X"d4019540",
		16#3c4e# => X"bd500007",
		16#3c4f# => X"0ffffef2",
		16#3c50# => X"d401853c",
		16#3c51# => X"03ffff0b",
		16#3c52# => X"84610028",
		16#3c53# => X"84610028",
		16#3c54# => X"84810020",
		16#3c55# => X"04001ac1",
		16#3c56# => X"9ca10538",
		16#3c57# => X"bc2b0000",
		16#3c58# => X"13fffb73",
		16#3c59# => X"9f0104d8",
		16#3c5a# => X"9ec104d0",
		16#3c5b# => X"86410540",
		16#3c5c# => X"03fffd5f",
		16#3c5d# => X"8601053c",
		16#3c5e# => X"0c0001e9",
		16#3c5f# => X"84410040",
		16#3c60# => X"9c600030",
		16#3c61# => X"9c42ffff",
		16#3c62# => X"d4011040",
		16#3c63# => X"d8021800",
		16#3c64# => X"84810014",
		16#3c65# => X"03fffbee",
		16#3c66# => X"e3441002",
		16#3c67# => X"e1c07002",
		16#3c68# => X"9c60002d",
		16#3c69# => X"e1607002",
		16#3c6a# => X"d8011d5b",
		16#3c6b# => X"e0eb7004",
		16#3c6c# => X"9d000001",
		16#3c6d# => X"03fffbc1",
		16#3c6e# => X"b967005f",
		16#3c6f# => X"9f050008",
		16#3c70# => X"8601053c",
		16#3c71# => X"aa948a3c",
		16#3c72# => X"9e100001",
		16#3c73# => X"e2527000",
		16#3c74# => X"d405a000",
		16#3c75# => X"d4057004",
		16#3c76# => X"d4019540",
		16#3c77# => X"bdb00007",
		16#3c78# => X"13fffd82",
		16#3c79# => X"d401853c",
		16#3c7a# => X"03fffe8b",
		16#3c7b# => X"84610028",
		16#3c7c# => X"85610050",
		16#3c7d# => X"a8ed0000",
		16#3c7e# => X"a90b0000",
		16#3c7f# => X"e0670004",
		16#3c80# => X"e0880004",
		16#3c81# => X"04001995",
		16#3c82# => X"15000000",
		16#3c83# => X"bc2b0000",
		16#3c84# => X"0c00015f",
		16#3c85# => X"18800001",
		16#3c86# => X"bc12ffff",
		16#3c87# => X"1000023e",
		16#3c88# => X"15000000",
		16#3c89# => X"ae1e0047",
		16#3c8a# => X"e1608002",
		16#3c8b# => X"e16b8004",
		16#3c8c# => X"bd6b0000",
		16#3c8d# => X"10000009",
		16#3c8e# => X"bc120000",
		16#3c8f# => X"ad9e0067",
		16#3c90# => X"e1606002",
		16#3c91# => X"e16b6004",
		16#3c92# => X"bd8b0000",
		16#3c93# => X"10000007",
		16#3c94# => X"84810018",
		16#3c95# => X"bc120000",
		16#3c96# => X"0c000004",
		16#3c97# => X"84810018",
		16#3c98# => X"9e400001",
		16#3c99# => X"84810018",
		16#3c9a# => X"8441004c",
		16#3c9b# => X"a8840100",
		16#3c9c# => X"bd620000",
		16#3c9d# => X"0c000224",
		16#3c9e# => X"d4012018",
		16#3c9f# => X"8701004c",
		16#3ca0# => X"9f800000",
		16#3ca1# => X"ac9e0046",
		16#3ca2# => X"ad7e0066",
		16#3ca3# => X"e0402002",
		16#3ca4# => X"e0605802",
		16#3ca5# => X"e0422004",
		16#3ca6# => X"e1635804",
		16#3ca7# => X"e16b1003",
		16#3ca8# => X"ad6bffff",
		16#3ca9# => X"bb4b005f",
		16#3caa# => X"bc3a0000",
		16#3cab# => X"100001fb",
		16#3cac# => X"a9d20000",
		16#3cad# => X"ad9e0045",
		16#3cae# => X"e1606002",
		16#3caf# => X"e16b6004",
		16#3cb0# => X"bd6b0000",
		16#3cb1# => X"10000009",
		16#3cb2# => X"9dd20001",
		16#3cb3# => X"ad9e0065",
		16#3cb4# => X"e1606002",
		16#3cb5# => X"e16b6004",
		16#3cb6# => X"bd8b0000",
		16#3cb7# => X"10000211",
		16#3cb8# => X"a9d20000",
		16#3cb9# => X"9dd20001",
		16#3cba# => X"9c400002",
		16#3cbb# => X"85e10050",
		16#3cbc# => X"a9980000",
		16#3cbd# => X"a9af0000",
		16#3cbe# => X"a8c20000",
		16#3cbf# => X"9c810550",
		16#3cc0# => X"84610028",
		16#3cc1# => X"a8ee0000",
		16#3cc2# => X"9d010554",
		16#3cc3# => X"9c41054c",
		16#3cc4# => X"d4012000",
		16#3cc5# => X"e08c0004",
		16#3cc6# => X"e0ad0004",
		16#3cc7# => X"04000491",
		16#3cc8# => X"d4011004",
		16#3cc9# => X"e1a08002",
		16#3cca# => X"e1ad8004",
		16#3ccb# => X"bd6d0000",
		16#3ccc# => X"10000008",
		16#3ccd# => X"d4015840",
		16#3cce# => X"ad9e0067",
		16#3ccf# => X"e1a06002",
		16#3cd0# => X"e1ad6004",
		16#3cd1# => X"bd8d0000",
		16#3cd2# => X"10000007",
		16#3cd3# => X"84810040",
		16#3cd4# => X"84610018",
		16#3cd5# => X"a5a30001",
		16#3cd6# => X"bc2d0000",
		16#3cd7# => X"0c0001f8",
		16#3cd8# => X"84810040",
		16#3cd9# => X"bc1a0000",
		16#3cda# => X"10000008",
		16#3cdb# => X"e0447000",
		16#3cdc# => X"91e40000",
		16#3cdd# => X"bc2f0030",
		16#3cde# => X"0c000202",
		16#3cdf# => X"85610050",
		16#3ce0# => X"85c10554",
		16#3ce1# => X"e0427000",
		16#3ce2# => X"84810050",
		16#3ce3# => X"18600001",
		16#3ce4# => X"a9980000",
		16#3ce5# => X"a86388d0",
		16#3ce6# => X"a9a40000",
		16#3ce7# => X"84a30000",
		16#3ce8# => X"84c30004",
		16#3ce9# => X"e06c0004",
		16#3cea# => X"e08d0004",
		16#3ceb# => X"07fff234",
		16#3cec# => X"15000000",
		16#3ced# => X"bc0b0000",
		16#3cee# => X"0c0001ba",
		16#3cef# => X"8461054c",
		16#3cf0# => X"d401154c",
		16#3cf1# => X"a8620000",
		16#3cf2# => X"84810040",
		16#3cf3# => X"e0408002",
		16#3cf4# => X"e0632002",
		16#3cf5# => X"e1028004",
		16#3cf6# => X"bd680000",
		16#3cf7# => X"10000008",
		16#3cf8# => X"d4011838",
		16#3cf9# => X"ad7e0067",
		16#3cfa# => X"e1005802",
		16#3cfb# => X"e1085804",
		16#3cfc# => X"bd880000",
		16#3cfd# => X"1000019a",
		16#3cfe# => X"bc1e0066",
		16#3cff# => X"87410554",
		16#3d00# => X"bd9afffd",
		16#3d01# => X"10000005",
		16#3d02# => X"a9da0000",
		16#3d03# => X"e572d000",
		16#3d04# => X"1000010c",
		16#3d05# => X"84810038",
		16#3d06# => X"9e9efffe",
		16#3d07# => X"9dceffff",
		16#3d08# => X"d801a544",
		16#3d09# => X"bd6e0000",
		16#3d0a# => X"0c0001cf",
		16#3d0b# => X"d4017554",
		16#3d0c# => X"9c60002b",
		16#3d0d# => X"d8011d45",
		16#3d0e# => X"bdae0009",
		16#3d0f# => X"100001bb",
		16#3d10# => X"9c800030",
		16#3d11# => X"9c41046f",
		16#3d12# => X"a86e0000",
		16#3d13# => X"9c80000a",
		16#3d14# => X"04002264",
		16#3d15# => X"9c42ffff",
		16#3d16# => X"9d6b0030",
		16#3d17# => X"a86e0000",
		16#3d18# => X"9c80000a",
		16#3d19# => X"07ffe8f2",
		16#3d1a# => X"d8025800",
		16#3d1b# => X"bd4b0009",
		16#3d1c# => X"13fffff6",
		16#3d1d# => X"a9cb0000",
		16#3d1e# => X"9d02ffff",
		16#3d1f# => X"9dcb0030",
		16#3d20# => X"d8087000",
		16#3d21# => X"8481000c",
		16#3d22# => X"e4682000",
		16#3d23# => X"10000009",
		16#3d24# => X"9ca10546",
		16#3d25# => X"8c480000",
		16#3d26# => X"d8051000",
		16#3d27# => X"9d080001",
		16#3d28# => X"8461000c",
		16#3d29# => X"e4881800",
		16#3d2a# => X"13fffffb",
		16#3d2b# => X"9ca50001",
		16#3d2c# => X"84410008",
		16#3d2d# => X"84610038",
		16#3d2e# => X"e0a51002",
		16#3d2f# => X"bd430001",
		16#3d30# => X"d4012858",
		16#3d31# => X"100000e7",
		16#3d32# => X"e3451800",
		16#3d33# => X"84810018",
		16#3d34# => X"a5040001",
		16#3d35# => X"bc080000",
		16#3d36# => X"0c0000e2",
		16#3d37# => X"15000000",
		16#3d38# => X"bc1c0000",
		16#3d39# => X"10000144",
		16#3d3a# => X"ac5affff",
		16#3d3b# => X"9c60002d",
		16#3d3c# => X"b842009f",
		16#3d3d# => X"9c800000",
		16#3d3e# => X"d8011d5b",
		16#3d3f# => X"e05a1003",
		16#3d40# => X"abd40000",
		16#3d41# => X"d4012044",
		16#3d42# => X"03fffb1a",
		16#3d43# => X"d4011024",
		16#3d44# => X"84610018",
		16#3d45# => X"a4430040",
		16#3d46# => X"bc020000",
		16#3d47# => X"10000096",
		16#3d48# => X"8481002c",
		16#3d49# => X"84610030",
		16#3d4a# => X"84440000",
		16#3d4b# => X"9c840004",
		16#3d4c# => X"d401202c",
		16#3d4d# => X"03fff9cb",
		16#3d4e# => X"dc021800",
		16#3d4f# => X"9d000001",
		16#3d50# => X"85c20000",
		16#3d51# => X"9c420004",
		16#3d52# => X"e1607002",
		16#3d53# => X"d401102c",
		16#3d54# => X"e0eb7004",
		16#3d55# => X"03fffbbc",
		16#3d56# => X"b967005f",
		16#3d57# => X"a90b0000",
		16#3d58# => X"85c30000",
		16#3d59# => X"9c630004",
		16#3d5a# => X"e1607002",
		16#3d5b# => X"d401182c",
		16#3d5c# => X"e0eb7004",
		16#3d5d# => X"03fffbb4",
		16#3d5e# => X"b967005f",
		16#3d5f# => X"a8b80000",
		16#3d60# => X"8601053c",
		16#3d61# => X"9f180008",
		16#3d62# => X"aa948a3c",
		16#3d63# => X"9e100001",
		16#3d64# => X"e2527000",
		16#3d65# => X"d405a000",
		16#3d66# => X"d4057004",
		16#3d67# => X"d4019540",
		16#3d68# => X"bdb00007",
		16#3d69# => X"1000000a",
		16#3d6a# => X"d401853c",
		16#3d6b# => X"84610028",
		16#3d6c# => X"84810020",
		16#3d6d# => X"040019a9",
		16#3d6e# => X"9ca10538",
		16#3d6f# => X"bc2b0000",
		16#3d70# => X"13fffa5b",
		16#3d71# => X"9f0104d0",
		16#3d72# => X"86410540",
		16#3d73# => X"84410018",
		16#3d74# => X"a4a20001",
		16#3d75# => X"bc050000",
		16#3d76# => X"13fffc85",
		16#3d77# => X"84810018",
		16#3d78# => X"8601053c",
		16#3d79# => X"84610054",
		16#3d7a# => X"9e100001",
		16#3d7b# => X"e2521800",
		16#3d7c# => X"84810048",
		16#3d7d# => X"d4182000",
		16#3d7e# => X"d4181804",
		16#3d7f# => X"d4019540",
		16#3d80# => X"bd500007",
		16#3d81# => X"13fffd83",
		16#3d82# => X"d401853c",
		16#3d83# => X"03fffc77",
		16#3d84# => X"9f180008",
		16#3d85# => X"1a800001",
		16#3d86# => X"a8b80000",
		16#3d87# => X"03fffc5b",
		16#3d88# => X"aa948a3c",
		16#3d89# => X"84610028",
		16#3d8a# => X"84810020",
		16#3d8b# => X"0400198b",
		16#3d8c# => X"9ca10538",
		16#3d8d# => X"bc2b0000",
		16#3d8e# => X"13fffa3d",
		16#3d8f# => X"9f0104d0",
		16#3d90# => X"03fffccf",
		16#3d91# => X"86410540",
		16#3d92# => X"19000001",
		16#3d93# => X"9e100001",
		16#3d94# => X"9e520001",
		16#3d95# => X"a908842b",
		16#3d96# => X"9c800001",
		16#3d97# => X"d4164000",
		16#3d98# => X"d4162004",
		16#3d99# => X"d4019540",
		16#3d9a# => X"bdb00007",
		16#3d9b# => X"0c000060",
		16#3d9c# => X"d401853c",
		16#3d9d# => X"bc2e0000",
		16#3d9e# => X"10000009",
		16#3d9f# => X"84410038",
		16#3da0# => X"bc220000",
		16#3da1# => X"10000006",
		16#3da2# => X"84610018",
		16#3da3# => X"a5030001",
		16#3da4# => X"bc080000",
		16#3da5# => X"13fffc56",
		16#3da6# => X"84810018",
		16#3da7# => X"8601053c",
		16#3da8# => X"84810054",
		16#3da9# => X"9e100001",
		16#3daa# => X"e2522000",
		16#3dab# => X"84410048",
		16#3dac# => X"d4182004",
		16#3dad# => X"d4181000",
		16#3dae# => X"d4019540",
		16#3daf# => X"bd500007",
		16#3db0# => X"10000055",
		16#3db1# => X"d401853c",
		16#3db2# => X"9f180008",
		16#3db3# => X"e1c07002",
		16#3db4# => X"bdae0000",
		16#3db5# => X"1000007c",
		16#3db6# => X"bdae0010",
		16#3db7# => X"10000094",
		16#3db8# => X"1a800001",
		16#3db9# => X"9c400010",
		16#3dba# => X"aa948a3c",
		16#3dbb# => X"86c10028",
		16#3dbc# => X"00000007",
		16#3dbd# => X"87410020",
		16#3dbe# => X"9f180008",
		16#3dbf# => X"9dcefff0",
		16#3dc0# => X"bd4e0010",
		16#3dc1# => X"0c00008b",
		16#3dc2# => X"15000000",
		16#3dc3# => X"9e100001",
		16#3dc4# => X"9e520010",
		16#3dc5# => X"d418a000",
		16#3dc6# => X"d4181004",
		16#3dc7# => X"d4019540",
		16#3dc8# => X"bd500007",
		16#3dc9# => X"0ffffff5",
		16#3dca# => X"d401853c",
		16#3dcb# => X"a8760000",
		16#3dcc# => X"a89a0000",
		16#3dcd# => X"04001949",
		16#3dce# => X"9ca10538",
		16#3dcf# => X"bc2b0000",
		16#3dd0# => X"13fff9fb",
		16#3dd1# => X"9f0104d0",
		16#3dd2# => X"86410540",
		16#3dd3# => X"03ffffec",
		16#3dd4# => X"8601053c",
		16#3dd5# => X"9c800000",
		16#3dd6# => X"b842009f",
		16#3dd7# => X"9101055b",
		16#3dd8# => X"e05a1003",
		16#3dd9# => X"d401702c",
		16#3dda# => X"d4012044",
		16#3ddb# => X"03fffa7e",
		16#3ddc# => X"d4011024",
		16#3ddd# => X"84610030",
		16#3dde# => X"84440000",
		16#3ddf# => X"9c840004",
		16#3de0# => X"d401202c",
		16#3de1# => X"03fff937",
		16#3de2# => X"d4021800",
		16#3de3# => X"bd5e0047",
		16#3de4# => X"a88488a2",
		16#3de5# => X"10000005",
		16#3de6# => X"d4012040",
		16#3de7# => X"18400001",
		16#3de8# => X"a842889e",
		16#3de9# => X"d4011040",
		16#3dea# => X"9c600003",
		16#3deb# => X"84810018",
		16#3dec# => X"9c40ff7f",
		16#3ded# => X"d4011824",
		16#3dee# => X"e0841003",
		16#3def# => X"ab430000",
		16#3df0# => X"9c600000",
		16#3df1# => X"d4012018",
		16#3df2# => X"9101055b",
		16#3df3# => X"03fffa66",
		16#3df4# => X"d4011844",
		16#3df5# => X"9d00002d",
		16#3df6# => X"03fffa90",
		16#3df7# => X"d8011d5b",
		16#3df8# => X"ab580000",
		16#3df9# => X"03fffd49",
		16#3dfa# => X"9f180008",
		16#3dfb# => X"84610028",
		16#3dfc# => X"84810020",
		16#3dfd# => X"04001919",
		16#3dfe# => X"9ca10538",
		16#3dff# => X"bc2b0000",
		16#3e00# => X"13fff9cb",
		16#3e01# => X"85c10554",
		16#3e02# => X"9f0104d0",
		16#3e03# => X"03ffff9a",
		16#3e04# => X"86410540",
		16#3e05# => X"84610028",
		16#3e06# => X"84810020",
		16#3e07# => X"0400190f",
		16#3e08# => X"9ca10538",
		16#3e09# => X"bc2b0000",
		16#3e0a# => X"13fff9c1",
		16#3e0b# => X"85c10554",
		16#3e0c# => X"9f0104d0",
		16#3e0d# => X"86410540",
		16#3e0e# => X"03ffffa5",
		16#3e0f# => X"8601053c",
		16#3e10# => X"e59a2000",
		16#3e11# => X"100000c0",
		16#3e12# => X"bd4e0000",
		16#3e13# => X"84610018",
		16#3e14# => X"a4430001",
		16#3e15# => X"bc020000",
		16#3e16# => X"13ffff22",
		16#3e17# => X"9e800067",
		16#3e18# => X"03ffff20",
		16#3e19# => X"9f5a0001",
		16#3e1a# => X"9f0e0008",
		16#3e1b# => X"03fffd27",
		16#3e1c# => X"ab4e0000",
		16#3e1d# => X"84610028",
		16#3e1e# => X"84810020",
		16#3e1f# => X"040018f7",
		16#3e20# => X"9ca10538",
		16#3e21# => X"bc2b0000",
		16#3e22# => X"13fff9a9",
		16#3e23# => X"86410540",
		16#3e24# => X"03fffc50",
		16#3e25# => X"9ca104d0",
		16#3e26# => X"03fffbd4",
		16#3e27# => X"ab050000",
		16#3e28# => X"84610028",
		16#3e29# => X"84810020",
		16#3e2a# => X"040018ec",
		16#3e2b# => X"9ca10538",
		16#3e2c# => X"bc2b0000",
		16#3e2d# => X"13fff99e",
		16#3e2e# => X"9f0104d0",
		16#3e2f# => X"86410540",
		16#3e30# => X"8601053c",
		16#3e31# => X"84610038",
		16#3e32# => X"9e100001",
		16#3e33# => X"e2521800",
		16#3e34# => X"03ffff49",
		16#3e35# => X"84810040",
		16#3e36# => X"07fff852",
		16#3e37# => X"d401702c",
		16#3e38# => X"adabffff",
		16#3e39# => X"9c400000",
		16#3e3a# => X"b9ad009f",
		16#3e3b# => X"ab4b0000",
		16#3e3c# => X"9101055b",
		16#3e3d# => X"e1ab6803",
		16#3e3e# => X"d4011044",
		16#3e3f# => X"03fffa1a",
		16#3e40# => X"d4016824",
		16#3e41# => X"1a800001",
		16#3e42# => X"9cf60008",
		16#3e43# => X"86410540",
		16#3e44# => X"8601053c",
		16#3e45# => X"03fff956",
		16#3e46# => X"aa948a4c",
		16#3e47# => X"84610014",
		16#3e48# => X"84810040",
		16#3e49# => X"03fffa0a",
		16#3e4a# => X"e3432002",
		16#3e4b# => X"aa948a3c",
		16#3e4c# => X"9e100001",
		16#3e4d# => X"e2527000",
		16#3e4e# => X"d418a000",
		16#3e4f# => X"d4187004",
		16#3e50# => X"d4019540",
		16#3e51# => X"bd500007",
		16#3e52# => X"13ffffd6",
		16#3e53# => X"d401853c",
		16#3e54# => X"03ffffdd",
		16#3e55# => X"9f180008",
		16#3e56# => X"bcb20006",
		16#3e57# => X"10000003",
		16#3e58# => X"ab520000",
		16#3e59# => X"9f400006",
		16#3e5a# => X"ac5affff",
		16#3e5b# => X"18800001",
		16#3e5c# => X"b842009f",
		16#3e5d# => X"a88488c8",
		16#3e5e# => X"d401702c",
		16#3e5f# => X"e05a1003",
		16#3e60# => X"d4012040",
		16#3e61# => X"03fff8fd",
		16#3e62# => X"d4011024",
		16#3e63# => X"84610028",
		16#3e64# => X"9c40ffff",
		16#3e65# => X"04000121",
		16#3e66# => X"d4011030",
		16#3e67# => X"bc2b0000",
		16#3e68# => X"13fff96b",
		16#3e69# => X"84610020",
		16#3e6a# => X"9843000c",
		16#3e6b# => X"03fff88f",
		16#3e6c# => X"a4e2ffff",
		16#3e6d# => X"1a800001",
		16#3e6e# => X"8601053c",
		16#3e6f# => X"03fffbb7",
		16#3e70# => X"aa948a4c",
		16#3e71# => X"84610028",
		16#3e72# => X"84810020",
		16#3e73# => X"040018a3",
		16#3e74# => X"9ca10538",
		16#3e75# => X"bc2b0000",
		16#3e76# => X"13fff955",
		16#3e77# => X"85c10554",
		16#3e78# => X"85610540",
		16#3e79# => X"a84e0000",
		16#3e7a# => X"8601053c",
		16#3e7b# => X"03fffc70",
		16#3e7c# => X"9f0104d0",
		16#3e7d# => X"9101055b",
		16#3e7e# => X"b842009f",
		16#3e7f# => X"abd40000",
		16#3e80# => X"d401e044",
		16#3e81# => X"e05a1003",
		16#3e82# => X"03fff9d7",
		16#3e83# => X"d4011024",
		16#3e84# => X"84610028",
		16#3e85# => X"84810020",
		16#3e86# => X"04001890",
		16#3e87# => X"9ca10538",
		16#3e88# => X"bc2b0000",
		16#3e89# => X"13fff942",
		16#3e8a# => X"85c10554",
		16#3e8b# => X"03fffc6b",
		16#3e8c# => X"9f0104d0",
		16#3e8d# => X"84610028",
		16#3e8e# => X"84810020",
		16#3e8f# => X"04001887",
		16#3e90# => X"9ca10538",
		16#3e91# => X"bc2b0000",
		16#3e92# => X"13fff939",
		16#3e93# => X"85c10554",
		16#3e94# => X"9f0104d0",
		16#3e95# => X"03fffd04",
		16#3e96# => X"86410540",
		16#3e97# => X"0c000046",
		16#3e98# => X"15000000",
		16#3e99# => X"87410554",
		16#3e9a# => X"bdba0000",
		16#3e9b# => X"1000005c",
		16#3e9c# => X"bc320000",
		16#3e9d# => X"10000006",
		16#3e9e# => X"84410018",
		16#3e9f# => X"a5020001",
		16#3ea0# => X"bc080000",
		16#3ea1# => X"13fffe98",
		16#3ea2# => X"bc1c0000",
		16#3ea3# => X"9f5a0001",
		16#3ea4# => X"03fffe94",
		16#3ea5# => X"e35a9000",
		16#3ea6# => X"03fffe15",
		16#3ea7# => X"9c400003",
		16#3ea8# => X"e4a21800",
		16#3ea9# => X"13fffe49",
		16#3eaa# => X"a8e30000",
		16#3eab# => X"9c800030",
		16#3eac# => X"d8072000",
		16#3ead# => X"9ce70001",
		16#3eae# => X"e4423800",
		16#3eaf# => X"13fffffd",
		16#3eb0# => X"d4013d4c",
		16#3eb1# => X"9da30001",
		16#3eb2# => X"9c800001",
		16#3eb3# => X"e1a46802",
		16#3eb4# => X"e1a26800",
		16#3eb5# => X"03fffe3d",
		16#3eb6# => X"e0636800",
		16#3eb7# => X"1a800001",
		16#3eb8# => X"a9180000",
		16#3eb9# => X"03fffc15",
		16#3eba# => X"aa948a3c",
		16#3ebb# => X"d4019024",
		16#3ebc# => X"9101055b",
		16#3ebd# => X"ab520000",
		16#3ebe# => X"d401702c",
		16#3ebf# => X"03fff99a",
		16#3ec0# => X"d4015844",
		16#3ec1# => X"18608000",
		16#3ec2# => X"9f80002d",
		16#3ec3# => X"03fffdde",
		16#3ec4# => X"e3021800",
		16#3ec5# => X"9e400006",
		16#3ec6# => X"03fffdd3",
		16#3ec7# => X"ae1e0047",
		16#3ec8# => X"03fffdf3",
		16#3ec9# => X"9c400002",
		16#3eca# => X"9dce0030",
		16#3ecb# => X"d8017547",
		16#3ecc# => X"d8012546",
		16#3ecd# => X"03fffe5f",
		16#3ece# => X"9ca10548",
		16#3ecf# => X"03fffe23",
		16#3ed0# => X"8461054c",
		16#3ed1# => X"10000004",
		16#3ed2# => X"9f400001",
		16#3ed3# => X"9c800002",
		16#3ed4# => X"e3447002",
		16#3ed5# => X"84410038",
		16#3ed6# => X"9e800067",
		16#3ed7# => X"03fffe61",
		16#3ed8# => X"e35a1000",
		16#3ed9# => X"9c40002d",
		16#3eda# => X"e1c07002",
		16#3edb# => X"03fffe33",
		16#3edc# => X"d8011545",
		16#3edd# => X"aa9e0000",
		16#3ede# => X"03fffe29",
		16#3edf# => X"85c10554",
		16#3ee0# => X"18600001",
		16#3ee1# => X"a9980000",
		16#3ee2# => X"a86388d0",
		16#3ee3# => X"a9ab0000",
		16#3ee4# => X"84a30000",
		16#3ee5# => X"84c30004",
		16#3ee6# => X"e06c0004",
		16#3ee7# => X"e08d0004",
		16#3ee8# => X"07fff055",
		16#3ee9# => X"15000000",
		16#3eea# => X"bc2b0000",
		16#3eeb# => X"0ffffdf5",
		16#3eec# => X"9c800001",
		16#3eed# => X"e1c47002",
		16#3eee# => X"03fffdf2",
		16#3eef# => X"d4017554",
		16#3ef0# => X"8441002c",
		16#3ef1# => X"86420000",
		16#3ef2# => X"bd920000",
		16#3ef3# => X"1000000f",
		16#3ef4# => X"9c420004",
		16#3ef5# => X"03fff857",
		16#3ef6# => X"d401102c",
		16#3ef7# => X"13fffe41",
		16#3ef8# => X"9f520002",
		16#3ef9# => X"84610018",
		16#3efa# => X"a4430001",
		16#3efb# => X"bc020000",
		16#3efc# => X"13fffe3c",
		16#3efd# => X"9f400001",
		16#3efe# => X"03fffe3a",
		16#3eff# => X"9f520002",
		16#3f00# => X"03fff905",
		16#3f01# => X"d4011830",
		16#3f02# => X"d401102c",
		16#3f03# => X"03fff849",
		16#3f04# => X"9e40ffff",
		16#3f05# => X"a8e40000",
		16#3f06# => X"a8830000",
		16#3f07# => X"18600001",
		16#3f08# => X"d7e14ffc",
		16#3f09# => X"a863ade4",
		16#3f0a# => X"9c21fffc",
		16#3f0b# => X"84630000",
		16#3f0c# => X"9c210004",
		16#3f0d# => X"a8c50000",
		16#3f0e# => X"8521fffc",
		16#3f0f# => X"03fff7b7",
		16#3f10# => X"a8a70000",
		16#3f11# => X"d7e117ec",
		16#3f12# => X"d7e187f4",
		16#3f13# => X"d7e197f8",
		16#3f14# => X"d7e14ffc",
		16#3f15# => X"d7e177f0",
		16#3f16# => X"aa030000",
		16#3f17# => X"9c21ffec",
		16#3f18# => X"aa440000",
		16#3f19# => X"bc030000",
		16#3f1a# => X"10000006",
		16#3f1b# => X"a8450000",
		16#3f1c# => X"84830038",
		16#3f1d# => X"bc240000",
		16#3f1e# => X"0c00003d",
		16#3f1f# => X"15000000",
		16#3f20# => X"98a2000c",
		16#3f21# => X"84820018",
		16#3f22# => X"a465ffff",
		16#3f23# => X"d4022008",
		16#3f24# => X"a4830008",
		16#3f25# => X"bc040000",
		16#3f26# => X"1000002b",
		16#3f27# => X"15000000",
		16#3f28# => X"84c20010",
		16#3f29# => X"bc260000",
		16#3f2a# => X"0c000027",
		16#3f2b# => X"15000000",
		16#3f2c# => X"a4632000",
		16#3f2d# => X"bc230000",
		16#3f2e# => X"0c00001d",
		16#3f2f# => X"9c80dfff",
		16#3f30# => X"84620000",
		16#3f31# => X"84820014",
		16#3f32# => X"e0c33002",
		16#3f33# => X"e5662000",
		16#3f34# => X"10000038",
		16#3f35# => X"9cc60001",
		16#3f36# => X"84a20008",
		16#3f37# => X"a5d200ff",
		16#3f38# => X"9ca5ffff",
		16#3f39# => X"9c830001",
		16#3f3a# => X"d4022808",
		16#3f3b# => X"d8037000",
		16#3f3c# => X"d4022000",
		16#3f3d# => X"84620014",
		16#3f3e# => X"e4033000",
		16#3f3f# => X"10000025",
		16#3f40# => X"bc2e000a",
		16#3f41# => X"0c00001e",
		16#3f42# => X"15000000",
		16#3f43# => X"9c210014",
		16#3f44# => X"a96e0000",
		16#3f45# => X"8521fffc",
		16#3f46# => X"8441ffec",
		16#3f47# => X"85c1fff0",
		16#3f48# => X"8601fff4",
		16#3f49# => X"44004800",
		16#3f4a# => X"8641fff8",
		16#3f4b# => X"84620064",
		16#3f4c# => X"a8a52000",
		16#3f4d# => X"e0632003",
		16#3f4e# => X"dc02280c",
		16#3f4f# => X"03ffffe1",
		16#3f50# => X"d4021864",
		16#3f51# => X"a8700000",
		16#3f52# => X"04000034",
		16#3f53# => X"a8820000",
		16#3f54# => X"bc2b0000",
		16#3f55# => X"10000020",
		16#3f56# => X"9dc0ffff",
		16#3f57# => X"98a2000c",
		16#3f58# => X"84c20010",
		16#3f59# => X"03ffffd3",
		16#3f5a# => X"a465ffff",
		16#3f5b# => X"04000a33",
		16#3f5c# => X"15000000",
		16#3f5d# => X"03ffffc4",
		16#3f5e# => X"98a2000c",
		16#3f5f# => X"9462000c",
		16#3f60# => X"a4630001",
		16#3f61# => X"bc030000",
		16#3f62# => X"13ffffe1",
		16#3f63# => X"15000000",
		16#3f64# => X"a8700000",
		16#3f65# => X"0400091b",
		16#3f66# => X"a8820000",
		16#3f67# => X"bc2b0000",
		16#3f68# => X"0fffffdb",
		16#3f69# => X"15000000",
		16#3f6a# => X"03ffffd9",
		16#3f6b# => X"9dc0ffff",
		16#3f6c# => X"a8700000",
		16#3f6d# => X"a8820000",
		16#3f6e# => X"04000912",
		16#3f6f# => X"9dc0ffff",
		16#3f70# => X"bc2b0000",
		16#3f71# => X"13ffffd2",
		16#3f72# => X"9cc00001",
		16#3f73# => X"03ffffc3",
		16#3f74# => X"84620000",
		16#3f75# => X"9462000c",
		16#3f76# => X"a8630040",
		16#3f77# => X"dc02180c",
		16#3f78# => X"9c400009",
		16#3f79# => X"03ffffca",
		16#3f7a# => X"d4101000",
		16#3f7b# => X"a8a40000",
		16#3f7c# => X"a8830000",
		16#3f7d# => X"18600001",
		16#3f7e# => X"d7e14ffc",
		16#3f7f# => X"a863ade4",
		16#3f80# => X"9c21fffc",
		16#3f81# => X"84630000",
		16#3f82# => X"9c210004",
		16#3f83# => X"8521fffc",
		16#3f84# => X"03ffff8d",
		16#3f85# => X"15000000",
		16#3f86# => X"d7e117f4",
		16#3f87# => X"18400001",
		16#3f88# => X"d7e177f8",
		16#3f89# => X"a842ade4",
		16#3f8a# => X"d7e14ffc",
		16#3f8b# => X"84a20000",
		16#3f8c# => X"9c21fff4",
		16#3f8d# => X"a9c30000",
		16#3f8e# => X"bc050000",
		16#3f8f# => X"10000006",
		16#3f90# => X"a8440000",
		16#3f91# => X"84650038",
		16#3f92# => X"bc230000",
		16#3f93# => X"0c00002b",
		16#3f94# => X"15000000",
		16#3f95# => X"98c2000c",
		16#3f96# => X"a486ffff",
		16#3f97# => X"a4640008",
		16#3f98# => X"bc030000",
		16#3f99# => X"10000032",
		16#3f9a# => X"a8e60000",
		16#3f9b# => X"84a20010",
		16#3f9c# => X"bc250000",
		16#3f9d# => X"0c000025",
		16#3f9e# => X"a4640280",
		16#3f9f# => X"a4640001",
		16#3fa0# => X"bc030000",
		16#3fa1# => X"1000000f",
		16#3fa2# => X"a4840002",
		16#3fa3# => X"84620014",
		16#3fa4# => X"9c800000",
		16#3fa5# => X"e0601802",
		16#3fa6# => X"9d600000",
		16#3fa7# => X"d4022008",
		16#3fa8# => X"e4255800",
		16#3fa9# => X"0c00000e",
		16#3faa# => X"d4021818",
		16#3fab# => X"9c21000c",
		16#3fac# => X"8521fffc",
		16#3fad# => X"8441fff4",
		16#3fae# => X"44004800",
		16#3faf# => X"85c1fff8",
		16#3fb0# => X"bc240000",
		16#3fb1# => X"10000003",
		16#3fb2# => X"9d600000",
		16#3fb3# => X"84620014",
		16#3fb4# => X"e4255800",
		16#3fb5# => X"13fffff6",
		16#3fb6# => X"d4021808",
		16#3fb7# => X"9442000c",
		16#3fb8# => X"a4420080",
		16#3fb9# => X"bc220000",
		16#3fba# => X"13fffff1",
		16#3fbb# => X"9d60ffff",
		16#3fbc# => X"03ffffef",
		16#3fbd# => X"a9650000",
		16#3fbe# => X"040009d0",
		16#3fbf# => X"a8650000",
		16#3fc0# => X"03ffffd6",
		16#3fc1# => X"98c2000c",
		16#3fc2# => X"bc030200",
		16#3fc3# => X"13ffffdd",
		16#3fc4# => X"a4640001",
		16#3fc5# => X"a8820000",
		16#3fc6# => X"04000dcb",
		16#3fc7# => X"a86e0000",
		16#3fc8# => X"9482000c",
		16#3fc9# => X"03ffffd6",
		16#3fca# => X"84a20010",
		16#3fcb# => X"a4640010",
		16#3fcc# => X"bc030000",
		16#3fcd# => X"13ffffde",
		16#3fce# => X"9d60ffff",
		16#3fcf# => X"a4840004",
		16#3fd0# => X"bc240000",
		16#3fd1# => X"10000007",
		16#3fd2# => X"15000000",
		16#3fd3# => X"84a20010",
		16#3fd4# => X"a8860008",
		16#3fd5# => X"dc02200c",
		16#3fd6# => X"03ffffc6",
		16#3fd7# => X"a484ffff",
		16#3fd8# => X"84820030",
		16#3fd9# => X"bc040000",
		16#3fda# => X"1000000a",
		16#3fdb# => X"9c620040",
		16#3fdc# => X"e4041800",
		16#3fdd# => X"10000006",
		16#3fde# => X"9c600000",
		16#3fdf# => X"04000ad0",
		16#3fe0# => X"a86e0000",
		16#3fe1# => X"98e2000c",
		16#3fe2# => X"9c600000",
		16#3fe3# => X"d4021830",
		16#3fe4# => X"84a20010",
		16#3fe5# => X"9c80ffdb",
		16#3fe6# => X"9c600000",
		16#3fe7# => X"e0c72003",
		16#3fe8# => X"d4021804",
		16#3fe9# => X"03ffffeb",
		16#3fea# => X"d4022800",
		16#3feb# => X"d7e117e4",
		16#3fec# => X"a8430000",
		16#3fed# => X"18600001",
		16#3fee# => X"d7e1b7f8",
		16#3fef# => X"a8638890",
		16#3ff0# => X"d7e187ec",
		16#3ff1# => X"86c30000",
		16#3ff2# => X"d7e197f0",
		16#3ff3# => X"d7e1a7f4",
		16#3ff4# => X"d7e14ffc",
		16#3ff5# => X"d7e177e8",
		16#3ff6# => X"84f60148",
		16#3ff7# => X"9c21ffe4",
		16#3ff8# => X"aa040000",
		16#3ff9# => X"aa850000",
		16#3ffa# => X"bc270000",
		16#3ffb# => X"0c00002c",
		16#3ffc# => X"aa460000",
		16#3ffd# => X"85070004",
		16#3ffe# => X"bda8001f",
		16#3fff# => X"0c00002b",
		16#4000# => X"18600000",
		16#4001# => X"bc020000",
		16#4002# => X"0c000013",
		16#4003# => X"9c880042",
		16#4004# => X"9c480002",
		16#4005# => X"9d080001",
		16#4006# => X"b8420002",
		16#4007# => X"d4074004",
		16#4008# => X"9dc00000",
		16#4009# => X"e0e71000",
		16#400a# => X"d4078000",
		16#400b# => X"9c21001c",
		16#400c# => X"a96e0000",
		16#400d# => X"8521fffc",
		16#400e# => X"8441ffe4",
		16#400f# => X"85c1ffe8",
		16#4010# => X"8601ffec",
		16#4011# => X"8641fff0",
		16#4012# => X"8681fff4",
		16#4013# => X"44004800",
		16#4014# => X"86c1fff8",
		16#4015# => X"9cc80022",
		16#4016# => X"9c600001",
		16#4017# => X"b8c60002",
		16#4018# => X"e0634008",
		16#4019# => X"b8840002",
		16#401a# => X"84a70188",
		16#401b# => X"e0c73000",
		16#401c# => X"e0a51804",
		16#401d# => X"e0872000",
		16#401e# => X"d406a000",
		16#401f# => X"d4072988",
		16#4020# => X"bc220002",
		16#4021# => X"13ffffe3",
		16#4022# => X"d4049000",
		16#4023# => X"8447018c",
		16#4024# => X"e0621804",
		16#4025# => X"03ffffdf",
		16#4026# => X"d407198c",
		16#4027# => X"9cf6014c",
		16#4028# => X"03ffffd5",
		16#4029# => X"d4163948",
		16#402a# => X"a863c5d8",
		16#402b# => X"bc030000",
		16#402c# => X"13ffffdf",
		16#402d# => X"9dc0ffff",
		16#402e# => X"07fff148",
		16#402f# => X"9c600190",
		16#4030# => X"bc0b0000",
		16#4031# => X"13ffffda",
		16#4032# => X"a8eb0000",
		16#4033# => X"84760148",
		16#4034# => X"9c800000",
		16#4035# => X"d40b1800",
		16#4036# => X"d40b2004",
		16#4037# => X"d4165948",
		16#4038# => X"d40b2188",
		16#4039# => X"d40b218c",
		16#403a# => X"03ffffc7",
		16#403b# => X"a9040000",
		16#403c# => X"d7e117d4",
		16#403d# => X"18400001",
		16#403e# => X"d7e1f7f8",
		16#403f# => X"a8428890",
		16#4040# => X"d7e1a7e4",
		16#4041# => X"87c20000",
		16#4042# => X"d7e1d7f0",
		16#4043# => X"d7e1e7f4",
		16#4044# => X"d7e14ffc",
		16#4045# => X"d7e177d8",
		16#4046# => X"d7e187dc",
		16#4047# => X"d7e197e0",
		16#4048# => X"d7e1b7e8",
		16#4049# => X"d7e1c7ec",
		16#404a# => X"9c5e0148",
		16#404b# => X"9c21ffd0",
		16#404c# => X"ab830000",
		16#404d# => X"aa840000",
		16#404e# => X"d4011000",
		16#404f# => X"9f400001",
		16#4050# => X"85de0148",
		16#4051# => X"bc0e0000",
		16#4052# => X"10000041",
		16#4053# => X"86c10000",
		16#4054# => X"848e0004",
		16#4055# => X"9c44ffff",
		16#4056# => X"bd820000",
		16#4057# => X"10000037",
		16#4058# => X"15000000",
		16#4059# => X"9e040021",
		16#405a# => X"9e440001",
		16#405b# => X"ba100002",
		16#405c# => X"ba520002",
		16#405d# => X"e20e8000",
		16#405e# => X"0000000b",
		16#405f# => X"e24e9000",
		16#4060# => X"84900080",
		16#4061# => X"e424a000",
		16#4062# => X"0c00000a",
		16#4063# => X"15000000",
		16#4064# => X"9c42ffff",
		16#4065# => X"9e10fffc",
		16#4066# => X"bd620000",
		16#4067# => X"0c000027",
		16#4068# => X"9e52fffc",
		16#4069# => X"bc140000",
		16#406a# => X"0ffffff6",
		16#406b# => X"15000000",
		16#406c# => X"848e0004",
		16#406d# => X"9c84ffff",
		16#406e# => X"e4241000",
		16#406f# => X"0c000035",
		16#4070# => X"84b20000",
		16#4071# => X"9c600000",
		16#4072# => X"d4121800",
		16#4073# => X"bc050000",
		16#4074# => X"13fffff0",
		16#4075# => X"e09a1008",
		16#4076# => X"84ce0188",
		16#4077# => X"e0c43003",
		16#4078# => X"bc260000",
		16#4079# => X"0c000027",
		16#407a# => X"870e0004",
		16#407b# => X"84ce018c",
		16#407c# => X"e0843003",
		16#407d# => X"bc240000",
		16#407e# => X"10000028",
		16#407f# => X"a87c0000",
		16#4080# => X"48002800",
		16#4081# => X"84900000",
		16#4082# => X"848e0004",
		16#4083# => X"e424c000",
		16#4084# => X"13ffffcc",
		16#4085# => X"15000000",
		16#4086# => X"84960000",
		16#4087# => X"e4247000",
		16#4088# => X"13ffffc8",
		16#4089# => X"9c42ffff",
		16#408a# => X"9e10fffc",
		16#408b# => X"bd620000",
		16#408c# => X"13ffffdd",
		16#408d# => X"9e52fffc",
		16#408e# => X"18400000",
		16#408f# => X"a842c600",
		16#4090# => X"bc020000",
		16#4091# => X"0c000019",
		16#4092# => X"15000000",
		16#4093# => X"9c210030",
		16#4094# => X"8521fffc",
		16#4095# => X"8441ffd4",
		16#4096# => X"85c1ffd8",
		16#4097# => X"8601ffdc",
		16#4098# => X"8641ffe0",
		16#4099# => X"8681ffe4",
		16#409a# => X"86c1ffe8",
		16#409b# => X"8701ffec",
		16#409c# => X"8741fff0",
		16#409d# => X"8781fff4",
		16#409e# => X"44004800",
		16#409f# => X"87c1fff8",
		16#40a0# => X"48002800",
		16#40a1# => X"15000000",
		16#40a2# => X"03ffffe1",
		16#40a3# => X"848e0004",
		16#40a4# => X"03ffffcf",
		16#40a5# => X"d40e1004",
		16#40a6# => X"48002800",
		16#40a7# => X"84700000",
		16#40a8# => X"03ffffdb",
		16#40a9# => X"848e0004",
		16#40aa# => X"844e0004",
		16#40ab# => X"bc220000",
		16#40ac# => X"0c00000a",
		16#40ad# => X"15000000",
		16#40ae# => X"844e0000",
		16#40af# => X"aace0000",
		16#40b0# => X"a9c20000",
		16#40b1# => X"bc2e0000",
		16#40b2# => X"13ffffa2",
		16#40b3# => X"15000000",
		16#40b4# => X"03ffffe0",
		16#40b5# => X"9c210030",
		16#40b6# => X"844e0000",
		16#40b7# => X"bc020000",
		16#40b8# => X"13fffff7",
		16#40b9# => X"a86e0000",
		16#40ba# => X"07fff0c6",
		16#40bb# => X"d4161000",
		16#40bc# => X"03fffff5",
		16#40bd# => X"85d60000",
		16#40be# => X"d7e117dc",
		16#40bf# => X"d7e177e0",
		16#40c0# => X"d7e187e4",
		16#40c1# => X"d7e1b7f0",
		16#40c2# => X"d7e1d7f8",
		16#40c3# => X"d7e14ffc",
		16#40c4# => X"d7e197e8",
		16#40c5# => X"d7e1a7ec",
		16#40c6# => X"d7e1c7f4",
		16#40c7# => X"84430010",
		16#40c8# => X"85c40010",
		16#40c9# => X"9c21ffdc",
		16#40ca# => X"aa030000",
		16#40cb# => X"aac40000",
		16#40cc# => X"e54e1000",
		16#40cd# => X"1000007f",
		16#40ce# => X"9f400000",
		16#40cf# => X"9c6e0004",
		16#40d0# => X"9c440014",
		16#40d1# => X"b8630002",
		16#40d2# => X"9dceffff",
		16#40d3# => X"9f100014",
		16#40d4# => X"e2441800",
		16#40d5# => X"e0701800",
		16#40d6# => X"84920000",
		16#40d7# => X"84630000",
		16#40d8# => X"07ffe4f4",
		16#40d9# => X"9c840001",
		16#40da# => X"e40bd000",
		16#40db# => X"1000003b",
		16#40dc# => X"aa8b0000",
		16#40dd# => X"a97a0000",
		16#40de# => X"a8c20000",
		16#40df# => X"a8b80000",
		16#40e0# => X"a87a0000",
		16#40e1# => X"85860000",
		16#40e2# => X"85050000",
		16#40e3# => X"a4ecffff",
		16#40e4# => X"b98c0050",
		16#40e5# => X"e0f43b06",
		16#40e6# => X"e1946306",
		16#40e7# => X"e0eb3800",
		16#40e8# => X"a488ffff",
		16#40e9# => X"b9670050",
		16#40ea# => X"e0632000",
		16#40eb# => X"a4e7ffff",
		16#40ec# => X"e16b6000",
		16#40ed# => X"e0833802",
		16#40ee# => X"b8680050",
		16#40ef# => X"a50bffff",
		16#40f0# => X"b8e40090",
		16#40f1# => X"e0634002",
		16#40f2# => X"a484ffff",
		16#40f3# => X"e0633800",
		16#40f4# => X"9cc60004",
		16#40f5# => X"b8e30010",
		16#40f6# => X"b96b0050",
		16#40f7# => X"b8630090",
		16#40f8# => X"e0872004",
		16#40f9# => X"e4723000",
		16#40fa# => X"d4052000",
		16#40fb# => X"13ffffe6",
		16#40fc# => X"9ca50004",
		16#40fd# => X"9cae0005",
		16#40fe# => X"b8a50002",
		16#40ff# => X"e0b02800",
		16#4100# => X"84650000",
		16#4101# => X"bc230000",
		16#4102# => X"10000015",
		16#4103# => X"a8700000",
		16#4104# => X"9ca5fffc",
		16#4105# => X"e4782800",
		16#4106# => X"1000000f",
		16#4107# => X"15000000",
		16#4108# => X"84650000",
		16#4109# => X"bc230000",
		16#410a# => X"0c000008",
		16#410b# => X"9ca5fffc",
		16#410c# => X"0000000a",
		16#410d# => X"d4107010",
		16#410e# => X"84650000",
		16#410f# => X"bc030000",
		16#4110# => X"0c000005",
		16#4111# => X"9ca5fffc",
		16#4112# => X"e4782800",
		16#4113# => X"0ffffffb",
		16#4114# => X"9dceffff",
		16#4115# => X"d4107010",
		16#4116# => X"a8700000",
		16#4117# => X"040010b4",
		16#4118# => X"a8960000",
		16#4119# => X"bd8b0000",
		16#411a# => X"10000031",
		16#411b# => X"a8980000",
		16#411c# => X"9e940001",
		16#411d# => X"9c600000",
		16#411e# => X"84e20000",
		16#411f# => X"85040000",
		16#4120# => X"a4a7ffff",
		16#4121# => X"a4c8ffff",
		16#4122# => X"b8e70050",
		16#4123# => X"e0a62802",
		16#4124# => X"b9080050",
		16#4125# => X"e0a51800",
		16#4126# => X"9c420004",
		16#4127# => X"b8c50090",
		16#4128# => X"e0683802",
		16#4129# => X"a4a5ffff",
		16#412a# => X"e0633000",
		16#412b# => X"e4721000",
		16#412c# => X"b8c30010",
		16#412d# => X"b8630090",
		16#412e# => X"e0a62804",
		16#412f# => X"d4042800",
		16#4130# => X"13ffffee",
		16#4131# => X"9c840004",
		16#4132# => X"9c4e0005",
		16#4133# => X"b8420002",
		16#4134# => X"e0501000",
		16#4135# => X"84620000",
		16#4136# => X"bc230000",
		16#4137# => X"10000015",
		16#4138# => X"ab540000",
		16#4139# => X"9c42fffc",
		16#413a# => X"e4781000",
		16#413b# => X"1000000f",
		16#413c# => X"15000000",
		16#413d# => X"84620000",
		16#413e# => X"bc230000",
		16#413f# => X"0c000008",
		16#4140# => X"9c42fffc",
		16#4141# => X"0000000b",
		16#4142# => X"d4107010",
		16#4143# => X"84620000",
		16#4144# => X"bc030000",
		16#4145# => X"0c000005",
		16#4146# => X"9c42fffc",
		16#4147# => X"e4781000",
		16#4148# => X"0ffffffb",
		16#4149# => X"9dceffff",
		16#414a# => X"d4107010",
		16#414b# => X"ab540000",
		16#414c# => X"9c210024",
		16#414d# => X"a97a0000",
		16#414e# => X"8521fffc",
		16#414f# => X"8441ffdc",
		16#4150# => X"85c1ffe0",
		16#4151# => X"8601ffe4",
		16#4152# => X"8641ffe8",
		16#4153# => X"8681ffec",
		16#4154# => X"86c1fff0",
		16#4155# => X"8701fff4",
		16#4156# => X"44004800",
		16#4157# => X"8741fff8",
		16#4158# => X"d7e117d4",
		16#4159# => X"d7e177d8",
		16#415a# => X"d7e1e7f4",
		16#415b# => X"d7e1f7f8",
		16#415c# => X"d7e14ffc",
		16#415d# => X"d7e187dc",
		16#415e# => X"d7e197e0",
		16#415f# => X"d7e1a7e4",
		16#4160# => X"d7e1b7e8",
		16#4161# => X"d7e1c7ec",
		16#4162# => X"d7e1d7f0",
		16#4163# => X"9c21ff64",
		16#4164# => X"84430040",
		16#4165# => X"d4013000",
		16#4166# => X"d4013818",
		16#4167# => X"d4014014",
		16#4168# => X"d4012810",
		16#4169# => X"abc30000",
		16#416a# => X"85c1009c",
		16#416b# => X"bc020000",
		16#416c# => X"1000000b",
		16#416d# => X"ab840000",
		16#416e# => X"85630044",
		16#416f# => X"9d800001",
		16#4170# => X"d4025804",
		16#4171# => X"e16c5808",
		16#4172# => X"a8820000",
		16#4173# => X"d4025808",
		16#4174# => X"04000e02",
		16#4175# => X"9c400000",
		16#4176# => X"d41e1040",
		16#4177# => X"bd7c0000",
		16#4178# => X"0c000204",
		16#4179# => X"9c800000",
		16#417a# => X"d40e2000",
		16#417b# => X"18c07ff0",
		16#417c# => X"e05c3003",
		16#417d# => X"e4223000",
		16#417e# => X"0c0001e2",
		16#417f# => X"85810010",
		16#4180# => X"18e00001",
		16#4181# => X"a85c0000",
		16#4182# => X"a86c0000",
		16#4183# => X"a8e78a6c",
		16#4184# => X"e0830004",
		16#4185# => X"e0620004",
		16#4186# => X"a9cc0000",
		16#4187# => X"84a70000",
		16#4188# => X"84c70004",
		16#4189# => X"07ffedb4",
		16#418a# => X"aa1c0000",
		16#418b# => X"bc2b0000",
		16#418c# => X"0c00001d",
		16#418d# => X"9c400001",
		16#418e# => X"a44200ff",
		16#418f# => X"bc220000",
		16#4190# => X"1000001f",
		16#4191# => X"ba5c0054",
		16#4192# => X"9c400001",
		16#4193# => X"84610014",
		16#4194# => X"19600001",
		16#4195# => X"848100a0",
		16#4196# => X"d4031000",
		16#4197# => X"bc040000",
		16#4198# => X"10000004",
		16#4199# => X"a96b842b",
		16#419a# => X"e04b1000",
		16#419b# => X"d4041000",
		16#419c# => X"9c21009c",
		16#419d# => X"8521fffc",
		16#419e# => X"8441ffd4",
		16#419f# => X"85c1ffd8",
		16#41a0# => X"8601ffdc",
		16#41a1# => X"8641ffe0",
		16#41a2# => X"8681ffe4",
		16#41a3# => X"86c1ffe8",
		16#41a4# => X"8701ffec",
		16#41a5# => X"8741fff0",
		16#41a6# => X"8781fff4",
		16#41a7# => X"44004800",
		16#41a8# => X"87c1fff8",
		16#41a9# => X"9c400000",
		16#41aa# => X"a44200ff",
		16#41ab# => X"bc220000",
		16#41ac# => X"0fffffe7",
		16#41ad# => X"9c400001",
		16#41ae# => X"ba5c0054",
		16#41af# => X"a9700000",
		16#41b0# => X"a98e0000",
		16#41b1# => X"a87e0000",
		16#41b2# => X"9cc10068",
		16#41b3# => X"9ce1006c",
		16#41b4# => X"e08b0004",
		16#41b5# => X"e0ac0004",
		16#41b6# => X"04001113",
		16#41b7# => X"a65207ff",
		16#41b8# => X"bc120000",
		16#41b9# => X"0c0001c9",
		16#41ba# => X"d4015830",
		16#41bb# => X"8681006c",
		16#41bc# => X"84410068",
		16#41bd# => X"e0541000",
		16#41be# => X"9e420432",
		16#41bf# => X"bdb20020",
		16#41c0# => X"10000368",
		16#41c1# => X"84810010",
		16#41c2# => X"9d800040",
		16#41c3# => X"9c420412",
		16#41c4# => X"e18c9002",
		16#41c5# => X"84610010",
		16#41c6# => X"e19c6008",
		16#41c7# => X"e0431048",
		16#41c8# => X"e04c1004",
		16#41c9# => X"a8620000",
		16#41ca# => X"07ffee5e",
		16#41cb# => X"9e52fbcd",
		16#41cc# => X"18c0fe10",
		16#41cd# => X"aa0b0000",
		16#41ce# => X"9ce00001",
		16#41cf# => X"e2103000",
		16#41d0# => X"a9cc0000",
		16#41d1# => X"d4013858",
		16#41d2# => X"a8500000",
		16#41d3# => X"a86e0000",
		16#41d4# => X"19800001",
		16#41d5# => X"e0830004",
		16#41d6# => X"e0620004",
		16#41d7# => X"18400001",
		16#41d8# => X"a98c8a74",
		16#41d9# => X"84ac0000",
		16#41da# => X"84cc0004",
		16#41db# => X"07ffeb0c",
		16#41dc# => X"a8428a7c",
		16#41dd# => X"84a20000",
		16#41de# => X"84c20004",
		16#41df# => X"18400001",
		16#41e0# => X"e06b0004",
		16#41e1# => X"e08c0004",
		16#41e2# => X"07ffeb27",
		16#41e3# => X"a8428a84",
		16#41e4# => X"84a20000",
		16#41e5# => X"84c20004",
		16#41e6# => X"e06b0004",
		16#41e7# => X"e08c0004",
		16#41e8# => X"07ffeae0",
		16#41e9# => X"18400001",
		16#41ea# => X"a8720000",
		16#41eb# => X"d4015808",
		16#41ec# => X"d401600c",
		16#41ed# => X"07ffee02",
		16#41ee# => X"a8428a8c",
		16#41ef# => X"84a20000",
		16#41f0# => X"84c20004",
		16#41f1# => X"e06b0004",
		16#41f2# => X"e08c0004",
		16#41f3# => X"07ffeb16",
		16#41f4# => X"15000000",
		16#41f5# => X"84610008",
		16#41f6# => X"8481000c",
		16#41f7# => X"e0ab0004",
		16#41f8# => X"e0cc0004",
		16#41f9# => X"07ffeacf",
		16#41fa# => X"15000000",
		16#41fb# => X"aa0b0000",
		16#41fc# => X"a86c0000",
		16#41fd# => X"a8500000",
		16#41fe# => X"e0830004",
		16#41ff# => X"e0620004",
		16#4200# => X"07ffee74",
		16#4201# => X"a9cc0000",
		16#4202# => X"18800001",
		16#4203# => X"a86e0000",
		16#4204# => X"a8848a6c",
		16#4205# => X"84a40000",
		16#4206# => X"84c40004",
		16#4207# => X"e0830004",
		16#4208# => X"e0620004",
		16#4209# => X"07ffed8e",
		16#420a# => X"d4015808",
		16#420b# => X"bd8b0000",
		16#420c# => X"0c000011",
		16#420d# => X"9ce00001",
		16#420e# => X"07ffede1",
		16#420f# => X"84610008",
		16#4210# => X"a9b00000",
		16#4211# => X"e06b0004",
		16#4212# => X"e08c0004",
		16#4213# => X"e0ad0004",
		16#4214# => X"e0ce0004",
		16#4215# => X"07ffed28",
		16#4216# => X"15000000",
		16#4217# => X"bc2b0000",
		16#4218# => X"0c000005",
		16#4219# => X"9ce00001",
		16#421a# => X"84c10008",
		16#421b# => X"9cc6ffff",
		16#421c# => X"d4013008",
		16#421d# => X"84410008",
		16#421e# => X"bc420016",
		16#421f# => X"10000017",
		16#4220# => X"d401383c",
		16#4221# => X"18600001",
		16#4222# => X"b9c20003",
		16#4223# => X"85e10010",
		16#4224# => X"a8638b04",
		16#4225# => X"a99c0000",
		16#4226# => X"a9af0000",
		16#4227# => X"e1ce1800",
		16#4228# => X"e0ac0004",
		16#4229# => X"e0cd0004",
		16#422a# => X"846e0000",
		16#422b# => X"848e0004",
		16#422c# => X"07ffed2f",
		16#422d# => X"15000000",
		16#422e# => X"bd4b0000",
		16#422f# => X"0c0002fd",
		16#4230# => X"9ce00000",
		16#4231# => X"84810008",
		16#4232# => X"9cc00000",
		16#4233# => X"9c84ffff",
		16#4234# => X"d401303c",
		16#4235# => X"d4012008",
		16#4236# => X"9e94ffff",
		16#4237# => X"e2549002",
		16#4238# => X"bd720000",
		16#4239# => X"0c0002ea",
		16#423a# => X"9c600000",
		16#423b# => X"d4019024",
		16#423c# => X"d4011834",
		16#423d# => X"84810008",
		16#423e# => X"bd840000",
		16#423f# => X"100002db",
		16#4240# => X"84c10024",
		16#4241# => X"9ce00000",
		16#4242# => X"e0c62000",
		16#4243# => X"d4012048",
		16#4244# => X"d4013024",
		16#4245# => X"d4013840",
		16#4246# => X"84e10000",
		16#4247# => X"bc470009",
		16#4248# => X"10000144",
		16#4249# => X"9c400000",
		16#424a# => X"bda70005",
		16#424b# => X"10000005",
		16#424c# => X"9dc00001",
		16#424d# => X"9ce7fffc",
		16#424e# => X"9dc00000",
		16#424f# => X"d4013800",
		16#4250# => X"84410000",
		16#4251# => X"bc020003",
		16#4252# => X"100004bc",
		16#4253# => X"bd420003",
		16#4254# => X"0c0002e8",
		16#4255# => X"bc020002",
		16#4256# => X"84610000",
		16#4257# => X"bc030004",
		16#4258# => X"100004b9",
		16#4259# => X"bc030005",
		16#425a# => X"0c0002e4",
		16#425b# => X"9cc0ffff",
		16#425c# => X"9c800001",
		16#425d# => X"d4012044",
		16#425e# => X"84c10008",
		16#425f# => X"84e10018",
		16#4260# => X"e0c63800",
		16#4261# => X"9e260001",
		16#4262# => X"bd510000",
		16#4263# => X"0c0004e3",
		16#4264# => X"d4013038",
		16#4265# => X"d401881c",
		16#4266# => X"9c400000",
		16#4267# => X"bc510017",
		16#4268# => X"0c00060b",
		16#4269# => X"d41e1044",
		16#426a# => X"9da00001",
		16#426b# => X"9d800004",
		16#426c# => X"e18c6000",
		16#426d# => X"a84d0000",
		16#426e# => X"9c6c0014",
		16#426f# => X"e4a38800",
		16#4270# => X"13fffffc",
		16#4271# => X"9dad0001",
		16#4272# => X"84c1001c",
		16#4273# => X"d41e1044",
		16#4274# => X"bca6000e",
		16#4275# => X"10000003",
		16#4276# => X"9d800001",
		16#4277# => X"9d800000",
		16#4278# => X"a87e0000",
		16#4279# => X"a8820000",
		16#427a# => X"04000ccf",
		16#427b# => X"e1ce6003",
		16#427c# => X"d4015820",
		16#427d# => X"bc0e0000",
		16#427e# => X"0c00011f",
		16#427f# => X"d41e5840",
		16#4280# => X"84c10008",
		16#4281# => X"85a10068",
		16#4282# => X"bda6000e",
		16#4283# => X"10000003",
		16#4284# => X"9d800001",
		16#4285# => X"9d800000",
		16#4286# => X"a58c00ff",
		16#4287# => X"bc0c0000",
		16#4288# => X"100001ee",
		16#4289# => X"84410044",
		16#428a# => X"bd8d0000",
		16#428b# => X"100001ec",
		16#428c# => X"bc020000",
		16#428d# => X"84e10008",
		16#428e# => X"18600001",
		16#428f# => X"b9870003",
		16#4290# => X"a8638b04",
		16#4291# => X"8441001c",
		16#4292# => X"e18c1800",
		16#4293# => X"bd420000",
		16#4294# => X"84cc0000",
		16#4295# => X"84ec0004",
		16#4296# => X"d4013000",
		16#4297# => X"d4013804",
		16#4298# => X"10000007",
		16#4299# => X"a9dc0000",
		16#429a# => X"84e10018",
		16#429b# => X"bd870000",
		16#429c# => X"10000353",
		16#429d# => X"84c1001c",
		16#429e# => X"a9dc0000",
		16#429f# => X"87810010",
		16#42a0# => X"84410020",
		16#42a1# => X"a8ee0000",
		16#42a2# => X"a91c0000",
		16#42a3# => X"9c420001",
		16#42a4# => X"e0670004",
		16#42a5# => X"e0880004",
		16#42a6# => X"84a10000",
		16#42a7# => X"84c10004",
		16#42a8# => X"07ffeb64",
		16#42a9# => X"d4011028",
		16#42aa# => X"e06b0004",
		16#42ab# => X"e08c0004",
		16#42ac# => X"07ffedc8",
		16#42ad# => X"15000000",
		16#42ae# => X"a86b0000",
		16#42af# => X"07ffed40",
		16#42b0# => X"aa4b0000",
		16#42b1# => X"84a10000",
		16#42b2# => X"84c10004",
		16#42b3# => X"e06b0004",
		16#42b4# => X"e08c0004",
		16#42b5# => X"07ffea54",
		16#42b6# => X"15000000",
		16#42b7# => X"a8ee0000",
		16#42b8# => X"a91c0000",
		16#42b9# => X"e0ab0004",
		16#42ba# => X"e0cc0004",
		16#42bb# => X"e0670004",
		16#42bc# => X"e0880004",
		16#42bd# => X"07ffea2a",
		16#42be# => X"15000000",
		16#42bf# => X"84610020",
		16#42c0# => X"a9ac0000",
		16#42c1# => X"9d920030",
		16#42c2# => X"a9cb0000",
		16#42c3# => X"d8036000",
		16#42c4# => X"a8ee0000",
		16#42c5# => X"8481001c",
		16#42c6# => X"bc040001",
		16#42c7# => X"1000005c",
		16#42c8# => X"a98d0000",
		16#42c9# => X"1b000001",
		16#42ca# => X"a8ee0000",
		16#42cb# => X"a90d0000",
		16#42cc# => X"ab188a9c",
		16#42cd# => X"e0670004",
		16#42ce# => X"e0880004",
		16#42cf# => X"84b80000",
		16#42d0# => X"84d80004",
		16#42d1# => X"07ffea38",
		16#42d2# => X"18400001",
		16#42d3# => X"a9cb0000",
		16#42d4# => X"a90c0000",
		16#42d5# => X"a8ee0000",
		16#42d6# => X"a8428a6c",
		16#42d7# => X"aa0c0000",
		16#42d8# => X"84a20000",
		16#42d9# => X"84c20004",
		16#42da# => X"e0670004",
		16#42db# => X"e0880004",
		16#42dc# => X"07ffec61",
		16#42dd# => X"9e400001",
		16#42de# => X"bc2b0000",
		16#42df# => X"10000004",
		16#42e0# => X"a65200ff",
		16#42e1# => X"aa4b0000",
		16#42e2# => X"a65200ff",
		16#42e3# => X"bc120000",
		16#42e4# => X"10000182",
		16#42e5# => X"9e800001",
		16#42e6# => X"8781001c",
		16#42e7# => X"00000017",
		16#42e8# => X"86c10028",
		16#42e9# => X"84b80000",
		16#42ea# => X"84d80004",
		16#42eb# => X"07ffea1e",
		16#42ec# => X"15000000",
		16#42ed# => X"18e00001",
		16#42ee# => X"a9cb0000",
		16#42ef# => X"a8e78a6c",
		16#42f0# => X"a86e0000",
		16#42f1# => X"a88c0000",
		16#42f2# => X"84a70000",
		16#42f3# => X"84c70004",
		16#42f4# => X"07ffec49",
		16#42f5# => X"aa0c0000",
		16#42f6# => X"bc2b0000",
		16#42f7# => X"10000004",
		16#42f8# => X"a75a00ff",
		16#42f9# => X"ab4b0000",
		16#42fa# => X"a75a00ff",
		16#42fb# => X"bc1a0000",
		16#42fc# => X"100004ce",
		16#42fd# => X"15000000",
		16#42fe# => X"a86e0000",
		16#42ff# => X"84a10000",
		16#4300# => X"84c10004",
		16#4301# => X"07ffeb0b",
		16#4302# => X"a8900000",
		16#4303# => X"e06b0004",
		16#4304# => X"e08c0004",
		16#4305# => X"07ffed6f",
		16#4306# => X"a84e0000",
		16#4307# => X"a86b0000",
		16#4308# => X"07ffece7",
		16#4309# => X"aa4b0000",
		16#430a# => X"84a10000",
		16#430b# => X"84c10004",
		16#430c# => X"e06b0004",
		16#430d# => X"e08c0004",
		16#430e# => X"07ffe9fb",
		16#430f# => X"9e940001",
		16#4310# => X"a8700000",
		16#4311# => X"e0ab0004",
		16#4312# => X"e0cc0004",
		16#4313# => X"e0830004",
		16#4314# => X"e0620004",
		16#4315# => X"07ffe9d2",
		16#4316# => X"9f400001",
		16#4317# => X"a88b0000",
		16#4318# => X"a8440000",
		16#4319# => X"9c920030",
		16#431a# => X"a86c0000",
		16#431b# => X"d8162000",
		16#431c# => X"e0830004",
		16#431d# => X"e0620004",
		16#431e# => X"e41ca000",
		16#431f# => X"0fffffca",
		16#4320# => X"9ed60001",
		16#4321# => X"d401b028",
		16#4322# => X"a8eb0000",
		16#4323# => X"a9a70000",
		16#4324# => X"a9cc0000",
		16#4325# => X"a8c70000",
		16#4326# => X"a8ec0000",
		16#4327# => X"e06d0004",
		16#4328# => X"e08e0004",
		16#4329# => X"e0a60004",
		16#432a# => X"e0c70004",
		16#432b# => X"07ffe99d",
		16#432c# => X"15000000",
		16#432d# => X"aa0b0000",
		16#432e# => X"a8ec0000",
		16#432f# => X"a8d00000",
		16#4330# => X"84410008",
		16#4331# => X"a9cc0000",
		16#4332# => X"84610000",
		16#4333# => X"84810004",
		16#4334# => X"e0a60004",
		16#4335# => X"e0c70004",
		16#4336# => X"07ffec61",
		16#4337# => X"d401105c",
		16#4338# => X"bd8b0000",
		16#4339# => X"10000013",
		16#433a# => X"84610028",
		16#433b# => X"a8ee0000",
		16#433c# => X"a8d00000",
		16#433d# => X"84610000",
		16#433e# => X"84810004",
		16#433f# => X"e0a60004",
		16#4340# => X"e0c70004",
		16#4341# => X"07ffebde",
		16#4342# => X"15000000",
		16#4343# => X"bc0b0000",
		16#4344# => X"0c000123",
		16#4345# => X"a87e0000",
		16#4346# => X"84610008",
		16#4347# => X"a6520001",
		16#4348# => X"bc320000",
		16#4349# => X"0c00011d",
		16#434a# => X"d401185c",
		16#434b# => X"84610028",
		16#434c# => X"00000003",
		16#434d# => X"84810020",
		16#434e# => X"a8620000",
		16#434f# => X"9c43ffff",
		16#4350# => X"90c20000",
		16#4351# => X"bc060039",
		16#4352# => X"0c000498",
		16#4353# => X"e4222000",
		16#4354# => X"13fffffa",
		16#4355# => X"9ce00030",
		16#4356# => X"d4012020",
		16#4357# => X"8481005c",
		16#4358# => X"84c10020",
		16#4359# => X"9c840001",
		16#435a# => X"d4011828",
		16#435b# => X"d4012008",
		16#435c# => X"d8063800",
		16#435d# => X"9cc00031",
		16#435e# => X"00000108",
		16#435f# => X"d8023000",
		16#4360# => X"9c40270f",
		16#4361# => X"84e10014",
		16#4362# => X"19600001",
		16#4363# => X"d4071000",
		16#4364# => X"84410010",
		16#4365# => X"bc220000",
		16#4366# => X"1000000b",
		16#4367# => X"a96b8a65",
		16#4368# => X"1860000f",
		16#4369# => X"19600001",
		16#436a# => X"a863ffff",
		16#436b# => X"e09c1803",
		16#436c# => X"bc040000",
		16#436d# => X"10000004",
		16#436e# => X"a96b8a5c",
		16#436f# => X"19600001",
		16#4370# => X"a96b8a65",
		16#4371# => X"848100a0",
		16#4372# => X"bc040000",
		16#4373# => X"13fffe29",
		16#4374# => X"9c4b0003",
		16#4375# => X"90620000",
		16#4376# => X"bc030000",
		16#4377# => X"10000003",
		16#4378# => X"84c100a0",
		16#4379# => X"9c4b0008",
		16#437a# => X"03fffe22",
		16#437b# => X"d4061000",
		16#437c# => X"18607fff",
		16#437d# => X"9c400001",
		16#437e# => X"a863ffff",
		16#437f# => X"d40e1000",
		16#4380# => X"03fffdfb",
		16#4381# => X"e39c1803",
		16#4382# => X"18c0000f",
		16#4383# => X"18e03ff0",
		16#4384# => X"a8c6ffff",
		16#4385# => X"9c400000",
		16#4386# => X"e2103003",
		16#4387# => X"9e52fc01",
		16#4388# => X"e2103804",
		16#4389# => X"8681006c",
		16#438a# => X"03fffe48",
		16#438b# => X"d4011058",
		16#438c# => X"9c60ffff",
		16#438d# => X"9c800001",
		16#438e# => X"d4011000",
		16#438f# => X"d4011838",
		16#4390# => X"a9c20000",
		16#4391# => X"d4012044",
		16#4392# => X"d401181c",
		16#4393# => X"d4011018",
		16#4394# => X"9c400000",
		16#4395# => X"d41e1044",
		16#4396# => X"a87e0000",
		16#4397# => X"04000bb2",
		16#4398# => X"a8820000",
		16#4399# => X"d4015820",
		16#439a# => X"bc0e0000",
		16#439b# => X"13fffee5",
		16#439c# => X"d41e5840",
		16#439d# => X"84e10010",
		16#439e# => X"84410008",
		16#439f# => X"d401382c",
		16#43a0# => X"bda20000",
		16#43a1# => X"100002b6",
		16#43a2# => X"aa5c0000",
		16#43a3# => X"a5e2000f",
		16#43a4# => X"18600001",
		16#43a5# => X"ba020084",
		16#43a6# => X"b9ef0003",
		16#43a7# => X"a8638b04",
		16#43a8# => X"a5d00010",
		16#43a9# => X"e1af1800",
		16#43aa# => X"9f400002",
		16#43ab# => X"bc0e0000",
		16#43ac# => X"86cd0000",
		16#43ad# => X"0c000181",
		16#43ae# => X"868d0004",
		16#43af# => X"bc100000",
		16#43b0# => X"10000014",
		16#43b1# => X"a9760000",
		16#43b2# => X"1b000001",
		16#43b3# => X"ab188bcc",
		16#43b4# => X"a9940000",
		16#43b5# => X"a4500001",
		16#43b6# => X"a86b0000",
		16#43b7# => X"a88c0000",
		16#43b8# => X"bc020000",
		16#43b9# => X"10000006",
		16#43ba# => X"ba100081",
		16#43bb# => X"84b80000",
		16#43bc# => X"84d80004",
		16#43bd# => X"07ffe94c",
		16#43be# => X"9f5a0001",
		16#43bf# => X"bc300000",
		16#43c0# => X"13fffff5",
		16#43c1# => X"9f180008",
		16#43c2# => X"aacb0000",
		16#43c3# => X"aa8c0000",
		16#43c4# => X"8581002c",
		16#43c5# => X"a8520000",
		16#43c6# => X"a9b60000",
		16#43c7# => X"a86c0000",
		16#43c8# => X"a9d40000",
		16#43c9# => X"e0830004",
		16#43ca# => X"e0620004",
		16#43cb# => X"e0ad0004",
		16#43cc# => X"e0ce0004",
		16#43cd# => X"07ffea3f",
		16#43ce# => X"15000000",
		16#43cf# => X"aa4b0000",
		16#43d0# => X"d401602c",
		16#43d1# => X"84e1003c",
		16#43d2# => X"bc070000",
		16#43d3# => X"1000003c",
		16#43d4# => X"a8520000",
		16#43d5# => X"85c1002c",
		16#43d6# => X"a86e0000",
		16#43d7# => X"19c00001",
		16#43d8# => X"e0830004",
		16#43d9# => X"e0620004",
		16#43da# => X"a9ce8a94",
		16#43db# => X"84ae0000",
		16#43dc# => X"84ce0004",
		16#43dd# => X"07ffebba",
		16#43de# => X"15000000",
		16#43df# => X"bd6b0000",
		16#43e0# => X"1000002f",
		16#43e1# => X"8441001c",
		16#43e2# => X"bda20000",
		16#43e3# => X"1000002c",
		16#43e4# => X"84610038",
		16#43e5# => X"bda30000",
		16#43e6# => X"13fffe9a",
		16#43e7# => X"8581002c",
		16#43e8# => X"1b000001",
		16#43e9# => X"a9b20000",
		16#43ea# => X"a9cc0000",
		16#43eb# => X"ab188a9c",
		16#43ec# => X"e06d0004",
		16#43ed# => X"e08e0004",
		16#43ee# => X"84b80000",
		16#43ef# => X"84d80004",
		16#43f0# => X"07ffe919",
		16#43f1# => X"1840fcc0",
		16#43f2# => X"84810008",
		16#43f3# => X"9c7a0001",
		16#43f4# => X"9c84ffff",
		16#43f5# => X"aa4b0000",
		16#43f6# => X"d401205c",
		16#43f7# => X"07ffebf8",
		16#43f8# => X"d401602c",
		16#43f9# => X"85a1002c",
		16#43fa# => X"84e10038",
		16#43fb# => X"a9ed0000",
		16#43fc# => X"a9d20000",
		16#43fd# => X"e0ab0004",
		16#43fe# => X"e0cc0004",
		16#43ff# => X"e06e0004",
		16#4400# => X"e08f0004",
		16#4401# => X"07ffe908",
		16#4402# => X"d401384c",
		16#4403# => X"1a600001",
		16#4404# => X"e06b0004",
		16#4405# => X"e08c0004",
		16#4406# => X"aa738aa4",
		16#4407# => X"84b30000",
		16#4408# => X"84d30004",
		16#4409# => X"07ffe8bf",
		16#440a# => X"15000000",
		16#440b# => X"aa8b0000",
		16#440c# => X"a9cc0000",
		16#440d# => X"00000140",
		16#440e# => X"e3541000",
		16#440f# => X"07ffebe0",
		16#4410# => X"a87a0000",
		16#4411# => X"85e1002c",
		16#4412# => X"a9b20000",
		16#4413# => X"a9cf0000",
		16#4414# => X"e06b0004",
		16#4415# => X"e08c0004",
		16#4416# => X"e0ad0004",
		16#4417# => X"e0ce0004",
		16#4418# => X"07ffe8f1",
		16#4419# => X"15000000",
		16#441a# => X"19a00001",
		16#441b# => X"e06b0004",
		16#441c# => X"e08c0004",
		16#441d# => X"a9ad8aa4",
		16#441e# => X"84ad0000",
		16#441f# => X"84cd0004",
		16#4420# => X"07ffe8a8",
		16#4421# => X"15000000",
		16#4422# => X"1860fcc0",
		16#4423# => X"a9ab0000",
		16#4424# => X"8481001c",
		16#4425# => X"ab0c0000",
		16#4426# => X"e34d1800",
		16#4427# => X"bc240000",
		16#4428# => X"10000121",
		16#4429# => X"a9cc0000",
		16#442a# => X"85e1002c",
		16#442b# => X"a8520000",
		16#442c# => X"a86f0000",
		16#442d# => X"19e00001",
		16#442e# => X"e0830004",
		16#442f# => X"e0620004",
		16#4430# => X"a9ef8aac",
		16#4431# => X"84af0000",
		16#4432# => X"84cf0004",
		16#4433# => X"07ffe8b4",
		16#4434# => X"aa180000",
		16#4435# => X"aacb0000",
		16#4436# => X"a9fa0000",
		16#4437# => X"aa760000",
		16#4438# => X"aa8c0000",
		16#4439# => X"e0730004",
		16#443a# => X"e0940004",
		16#443b# => X"e0af0004",
		16#443c# => X"e0d00004",
		16#443d# => X"07ffeb1e",
		16#443e# => X"a9cc0000",
		16#443f# => X"bd4b0000",
		16#4440# => X"100001c5",
		16#4441# => X"18c08000",
		16#4442# => X"a9f60000",
		16#4443# => X"e2ba3000",
		16#4444# => X"aa0e0000",
		16#4445# => X"a9b50000",
		16#4446# => X"a9d80000",
		16#4447# => X"e06f0004",
		16#4448# => X"e0900004",
		16#4449# => X"e0ad0004",
		16#444a# => X"e0ce0004",
		16#444b# => X"07ffeb4c",
		16#444c# => X"15000000",
		16#444d# => X"bd8b0000",
		16#444e# => X"0ffffe33",
		16#444f# => X"84c10008",
		16#4450# => X"8441001c",
		16#4451# => X"aa420000",
		16#4452# => X"84810018",
		16#4453# => X"84c10020",
		16#4454# => X"ac84ffff",
		16#4455# => X"d4013028",
		16#4456# => X"d4012008",
		16#4457# => X"9dc00000",
		16#4458# => X"a87e0000",
		16#4459# => X"04000b1d",
		16#445a# => X"a8820000",
		16#445b# => X"bc120000",
		16#445c# => X"1000000a",
		16#445d# => X"e0ce9005",
		16#445e# => X"e0e03002",
		16#445f# => X"e0c73004",
		16#4460# => X"bd660000",
		16#4461# => X"0c0001e2",
		16#4462# => X"e0c07002",
		16#4463# => X"a87e0000",
		16#4464# => X"04000b12",
		16#4465# => X"a8920000",
		16#4466# => X"a87e0000",
		16#4467# => X"04000b0f",
		16#4468# => X"84810030",
		16#4469# => X"84610028",
		16#446a# => X"9c800000",
		16#446b# => X"84e10008",
		16#446c# => X"d8032000",
		16#446d# => X"9c470001",
		16#446e# => X"84c10014",
		16#446f# => X"84e100a0",
		16#4470# => X"d4061000",
		16#4471# => X"bc070000",
		16#4472# => X"13fffd2a",
		16#4473# => X"85610020",
		16#4474# => X"03fffd28",
		16#4475# => X"d4071800",
		16#4476# => X"bc020000",
		16#4477# => X"100000ce",
		16#4478# => X"84610000",
		16#4479# => X"bd430001",
		16#447a# => X"0c000368",
		16#447b# => X"84c1001c",
		16#447c# => X"84e10040",
		16#447d# => X"9e06ffff",
		16#447e# => X"e5878000",
		16#447f# => X"10000353",
		16#4480# => X"84410040",
		16#4481# => X"e2078002",
		16#4482# => X"8481001c",
		16#4483# => X"bd640000",
		16#4484# => X"0c000375",
		16#4485# => X"84c10034",
		16#4486# => X"85c10034",
		16#4487# => X"85a1001c",
		16#4488# => X"84e10034",
		16#4489# => X"84410024",
		16#448a# => X"e0e76800",
		16#448b# => X"e0426800",
		16#448c# => X"a87e0000",
		16#448d# => X"9c800001",
		16#448e# => X"d4013834",
		16#448f# => X"04000be7",
		16#4490# => X"d4011024",
		16#4491# => X"aa4b0000",
		16#4492# => X"84610024",
		16#4493# => X"bda30000",
		16#4494# => X"1000000f",
		16#4495# => X"bdae0000",
		16#4496# => X"1000000e",
		16#4497# => X"84e10040",
		16#4498# => X"e5a37000",
		16#4499# => X"10000003",
		16#449a# => X"a9830000",
		16#449b# => X"a98e0000",
		16#449c# => X"84810034",
		16#449d# => X"84c10024",
		16#449e# => X"e0846002",
		16#449f# => X"e0c66002",
		16#44a0# => X"d4012034",
		16#44a1# => X"e1ce6002",
		16#44a2# => X"d4013024",
		16#44a3# => X"84e10040",
		16#44a4# => X"bda70000",
		16#44a5# => X"10000018",
		16#44a6# => X"84410044",
		16#44a7# => X"bc020000",
		16#44a8# => X"10000324",
		16#44a9# => X"bdb00000",
		16#44aa# => X"1000000e",
		16#44ab# => X"a8920000",
		16#44ac# => X"a87e0000",
		16#44ad# => X"04000c67",
		16#44ae# => X"a8b00000",
		16#44af# => X"a87e0000",
		16#44b0# => X"a88b0000",
		16#44b1# => X"84a10030",
		16#44b2# => X"04000bd1",
		16#44b3# => X"aa4b0000",
		16#44b4# => X"84810030",
		16#44b5# => X"a87e0000",
		16#44b6# => X"04000ac0",
		16#44b7# => X"d4015830",
		16#44b8# => X"84610040",
		16#44b9# => X"e2038002",
		16#44ba# => X"bc100000",
		16#44bb# => X"0c00031f",
		16#44bc# => X"a87e0000",
		16#44bd# => X"9c800001",
		16#44be# => X"04000bb8",
		16#44bf# => X"a87e0000",
		16#44c0# => X"84810048",
		16#44c1# => X"bda40000",
		16#44c2# => X"10000007",
		16#44c3# => X"a84b0000",
		16#44c4# => X"a87e0000",
		16#44c5# => X"a88b0000",
		16#44c6# => X"04000c4e",
		16#44c7# => X"84a10048",
		16#44c8# => X"a84b0000",
		16#44c9# => X"84c10000",
		16#44ca# => X"bd460001",
		16#44cb# => X"0c000282",
		16#44cc# => X"9e000000",
		16#44cd# => X"84610048",
		16#44ce# => X"bc030000",
		16#44cf# => X"0c000269",
		16#44d0# => X"9da00001",
		16#44d1# => X"84810024",
		16#44d2# => X"e1ad2000",
		16#44d3# => X"a5ad001f",
		16#44d4# => X"bc0d0000",
		16#44d5# => X"0c000176",
		16#44d6# => X"9d80001c",
		16#44d7# => X"84e10034",
		16#44d8# => X"84610024",
		16#44d9# => X"e0e76000",
		16#44da# => X"e0636000",
		16#44db# => X"d4013834",
		16#44dc# => X"e1ce6000",
		16#44dd# => X"d4011824",
		16#44de# => X"84810034",
		16#44df# => X"bda40000",
		16#44e0# => X"10000008",
		16#44e1# => X"84c10024",
		16#44e2# => X"a87e0000",
		16#44e3# => X"84810030",
		16#44e4# => X"04000c88",
		16#44e5# => X"84a10034",
		16#44e6# => X"d4015830",
		16#44e7# => X"84c10024",
		16#44e8# => X"bda60000",
		16#44e9# => X"10000008",
		16#44ea# => X"84e1003c",
		16#44eb# => X"a8820000",
		16#44ec# => X"a87e0000",
		16#44ed# => X"04000c7f",
		16#44ee# => X"a8a60000",
		16#44ef# => X"a84b0000",
		16#44f0# => X"84e1003c",
		16#44f1# => X"bc070000",
		16#44f2# => X"0c00022b",
		16#44f3# => X"15000000",
		16#44f4# => X"84c1001c",
		16#44f5# => X"bd460000",
		16#44f6# => X"10000112",
		16#44f7# => X"84e10044",
		16#44f8# => X"84e10000",
		16#44f9# => X"bd470002",
		16#44fa# => X"10000003",
		16#44fb# => X"9d800001",
		16#44fc# => X"9d800000",
		16#44fd# => X"a58c00ff",
		16#44fe# => X"bc0c0000",
		16#44ff# => X"10000109",
		16#4500# => X"84e10044",
		16#4501# => X"8461001c",
		16#4502# => X"bc230000",
		16#4503# => X"13ffff4f",
		16#4504# => X"a8c30000",
		16#4505# => X"a8820000",
		16#4506# => X"9ca00005",
		16#4507# => X"04000a7b",
		16#4508# => X"a87e0000",
		16#4509# => X"84610030",
		16#450a# => X"a88b0000",
		16#450b# => X"04000cc0",
		16#450c# => X"a84b0000",
		16#450d# => X"bd4b0000",
		16#450e# => X"0fffff44",
		16#450f# => X"15000000",
		16#4510# => X"84e10020",
		16#4511# => X"9c600031",
		16#4512# => X"9c870001",
		16#4513# => X"d8071800",
		16#4514# => X"d4012028",
		16#4515# => X"84c10008",
		16#4516# => X"9dc00000",
		16#4517# => X"9cc60001",
		16#4518# => X"03ffff40",
		16#4519# => X"d4013008",
		16#451a# => X"84410034",
		16#451b# => X"84610008",
		16#451c# => X"9cc00000",
		16#451d# => X"e0421802",
		16#451e# => X"e0801802",
		16#451f# => X"d4011034",
		16#4520# => X"d4012040",
		16#4521# => X"03fffd25",
		16#4522# => X"d4013048",
		16#4523# => X"e2409002",
		16#4524# => X"9c400000",
		16#4525# => X"d4019034",
		16#4526# => X"03fffd17",
		16#4527# => X"d4011024",
		16#4528# => X"9c400020",
		16#4529# => X"e0429002",
		16#452a# => X"03fffc9f",
		16#452b# => X"e0441008",
		16#452c# => X"03fffd0a",
		16#452d# => X"d401383c",
		16#452e# => X"19800001",
		16#452f# => X"a8670000",
		16#4530# => X"a98c8bcc",
		16#4531# => X"a85c0000",
		16#4532# => X"84ac0020",
		16#4533# => X"84cc0024",
		16#4534# => X"e0830004",
		16#4535# => X"e0620004",
		16#4536# => X"07ffe8d6",
		16#4537# => X"a610000f",
		16#4538# => X"9f400003",
		16#4539# => X"aa4b0000",
		16#453a# => X"03fffe75",
		16#453b# => X"d401602c",
		16#453c# => X"100001de",
		16#453d# => X"9cc0ffff",
		16#453e# => X"9dc00000",
		16#453f# => X"9ce00001",
		16#4540# => X"d4013038",
		16#4541# => X"d4013844",
		16#4542# => X"d401301c",
		16#4543# => X"03fffe51",
		16#4544# => X"d4017018",
		16#4545# => X"86010040",
		16#4546# => X"85c10034",
		16#4547# => X"03ffff4b",
		16#4548# => X"86410044",
		16#4549# => X"84e10008",
		16#454a# => X"8441001c",
		16#454b# => X"d401385c",
		16#454c# => X"d401104c",
		16#454d# => X"84610044",
		16#454e# => X"bc030000",
		16#454f# => X"10000136",
		16#4550# => X"8481004c",
		16#4551# => X"18c00001",
		16#4552# => X"9e64ffff",
		16#4553# => X"a8c68b04",
		16#4554# => X"ba730003",
		16#4555# => X"e1933000",
		16#4556# => X"1a600001",
		16#4557# => X"84ac0000",
		16#4558# => X"84cc0004",
		16#4559# => X"aa738ab4",
		16#455a# => X"84730000",
		16#455b# => X"84930004",
		16#455c# => X"07ffe8b0",
		16#455d# => X"aada0000",
		16#455e# => X"84e10020",
		16#455f# => X"aaee0000",
		16#4560# => X"9ce70001",
		16#4561# => X"e0b60004",
		16#4562# => X"e0d70004",
		16#4563# => X"e06b0004",
		16#4564# => X"e08c0004",
		16#4565# => X"07ffe782",
		16#4566# => X"d4013828",
		16#4567# => X"8461002c",
		16#4568# => X"aab20000",
		16#4569# => X"aac30000",
		16#456a# => X"aa0c0000",
		16#456b# => X"e0750004",
		16#456c# => X"e0960004",
		16#456d# => X"07ffeb07",
		16#456e# => X"aa8b0000",
		16#456f# => X"a86b0000",
		16#4570# => X"07ffea7f",
		16#4571# => X"a84b0000",
		16#4572# => X"85e1002c",
		16#4573# => X"aab20000",
		16#4574# => X"aacf0000",
		16#4575# => X"e0ab0004",
		16#4576# => X"e0cc0004",
		16#4577# => X"e0750004",
		16#4578# => X"e0960004",
		16#4579# => X"07ffe76e",
		16#457a# => X"aad00000",
		16#457b# => X"9ce20030",
		16#457c# => X"ab4b0000",
		16#457d# => X"84410020",
		16#457e# => X"aab40000",
		16#457f# => X"a9ba0000",
		16#4580# => X"a9cc0000",
		16#4581# => X"d8023800",
		16#4582# => X"e0750004",
		16#4583# => X"e0960004",
		16#4584# => X"e0ad0004",
		16#4585# => X"e0ce0004",
		16#4586# => X"07ffe9d5",
		16#4587# => X"aa4c0000",
		16#4588# => X"bd4b0000",
		16#4589# => X"100002e7",
		16#458a# => X"18c00001",
		16#458b# => X"a9ba0000",
		16#458c# => X"a8c68a94",
		16#458d# => X"84660000",
		16#458e# => X"84860004",
		16#458f# => X"e0ad0004",
		16#4590# => X"e0ce0004",
		16#4591# => X"07ffe756",
		16#4592# => X"a9d00000",
		16#4593# => X"a9b40000",
		16#4594# => X"e0ab0004",
		16#4595# => X"e0cc0004",
		16#4596# => X"e06d0004",
		16#4597# => X"e08e0004",
		16#4598# => X"07ffe9c3",
		16#4599# => X"15000000",
		16#459a# => X"bd4b0000",
		16#459b# => X"13fffdb0",
		16#459c# => X"84e1004c",
		16#459d# => X"bda70001",
		16#459e# => X"13fffce2",
		16#459f# => X"1b000001",
		16#45a0# => X"9ec00001",
		16#45a1# => X"ab188a9c",
		16#45a2# => X"d401f060",
		16#45a3# => X"85d80000",
		16#45a4# => X"87180004",
		16#45a5# => X"d401e064",
		16#45a6# => X"d401c050",
		16#45a7# => X"ab960000",
		16#45a8# => X"d401c054",
		16#45a9# => X"d401702c",
		16#45aa# => X"aad00000",
		16#45ab# => X"abce0000",
		16#45ac# => X"00000014",
		16#45ad# => X"87010028",
		16#45ae# => X"18400001",
		16#45af# => X"a8428a94",
		16#45b0# => X"84620000",
		16#45b1# => X"84820004",
		16#45b2# => X"07ffe735",
		16#45b3# => X"15000000",
		16#45b4# => X"a8b40000",
		16#45b5# => X"e06b0004",
		16#45b6# => X"e08c0004",
		16#45b7# => X"07ffe9e0",
		16#45b8# => X"a8d60000",
		16#45b9# => X"bd8b0000",
		16#45ba# => X"10000239",
		16#45bb# => X"a8780000",
		16#45bc# => X"8461004c",
		16#45bd# => X"e57c1800",
		16#45be# => X"10000238",
		16#45bf# => X"15000000",
		16#45c0# => X"a8740000",
		16#45c1# => X"a8960000",
		16#45c2# => X"84c10054",
		16#45c3# => X"a8be0000",
		16#45c4# => X"07ffe745",
		16#45c5# => X"9f9c0001",
		16#45c6# => X"84a1002c",
		16#45c7# => X"84c10050",
		16#45c8# => X"a87a0000",
		16#45c9# => X"a8920000",
		16#45ca# => X"aa8b0000",
		16#45cb# => X"07ffe73e",
		16#45cc# => X"aacc0000",
		16#45cd# => X"aa4b0000",
		16#45ce# => X"a88c0000",
		16#45cf# => X"a8720000",
		16#45d0# => X"07ffeaa4",
		16#45d1# => X"aa0c0000",
		16#45d2# => X"a86b0000",
		16#45d3# => X"07ffea1c",
		16#45d4# => X"a9cb0000",
		16#45d5# => X"a8520000",
		16#45d6# => X"a8700000",
		16#45d7# => X"e0ab0004",
		16#45d8# => X"e0cc0004",
		16#45d9# => X"e0830004",
		16#45da# => X"e0620004",
		16#45db# => X"07ffe70c",
		16#45dc# => X"9dce0030",
		16#45dd# => X"ab4b0000",
		16#45de# => X"a8b40000",
		16#45df# => X"d8187000",
		16#45e0# => X"a8d60000",
		16#45e1# => X"a87a0000",
		16#45e2# => X"a88c0000",
		16#45e3# => X"07ffe9b4",
		16#45e4# => X"aa4c0000",
		16#45e5# => X"9f180001",
		16#45e6# => X"a8ba0000",
		16#45e7# => X"bd8b0000",
		16#45e8# => X"0fffffc6",
		16#45e9# => X"a8d20000",
		16#45ea# => X"84c1005c",
		16#45eb# => X"d401c028",
		16#45ec# => X"87c10060",
		16#45ed# => X"03fffe79",
		16#45ee# => X"d4013008",
		16#45ef# => X"bc260000",
		16#45f0# => X"100001ef",
		16#45f1# => X"19800001",
		16#45f2# => X"84610000",
		16#45f3# => X"84810004",
		16#45f4# => X"a98c8aac",
		16#45f5# => X"84ac0000",
		16#45f6# => X"84cc0004",
		16#45f7# => X"07ffe712",
		16#45f8# => X"a9dc0000",
		16#45f9# => X"87810010",
		16#45fa# => X"e06b0004",
		16#45fb# => X"e08c0004",
		16#45fc# => X"a9bc0000",
		16#45fd# => X"a98e0000",
		16#45fe# => X"e0ac0004",
		16#45ff# => X"e0cd0004",
		16#4600# => X"07ffe979",
		16#4601# => X"15000000",
		16#4602# => X"bd6b0000",
		16#4603# => X"13fffe4d",
		16#4604# => X"15000000",
		16#4605# => X"8441001c",
		16#4606# => X"03ffff0a",
		16#4607# => X"aa420000",
		16#4608# => X"bc270000",
		16#4609# => X"1000015b",
		16#460a# => X"bdae0000",
		16#460b# => X"84610020",
		16#460c# => X"9dc00001",
		16#460d# => X"d4011828",
		16#460e# => X"8601001c",
		16#460f# => X"86c10030",
		16#4610# => X"00000005",
		16#4611# => X"aa830000",
		16#4612# => X"04000970",
		16#4613# => X"9dce0001",
		16#4614# => X"aacb0000",
		16#4615# => X"a8760000",
		16#4616# => X"07fffaa8",
		16#4617# => X"a8820000",
		16#4618# => X"9d6b0030",
		16#4619# => X"a87e0000",
		16#461a# => X"d8145800",
		16#461b# => X"a8960000",
		16#461c# => X"9ca0000a",
		16#461d# => X"9cc00000",
		16#461e# => X"e56e8000",
		16#461f# => X"0ffffff3",
		16#4620# => X"9e940001",
		16#4621# => X"aa0b0000",
		16#4622# => X"d401b030",
		16#4623# => X"d401a028",
		16#4624# => X"9dc00000",
		16#4625# => X"9ca00001",
		16#4626# => X"a87e0000",
		16#4627# => X"04000b45",
		16#4628# => X"84810030",
		16#4629# => X"a8820000",
		16#462a# => X"a86b0000",
		16#462b# => X"04000ba0",
		16#462c# => X"d4015830",
		16#462d# => X"bd4b0000",
		16#462e# => X"0c0001e6",
		16#462f# => X"bc2b0000",
		16#4630# => X"84610028",
		16#4631# => X"00000003",
		16#4632# => X"84810020",
		16#4633# => X"a8660000",
		16#4634# => X"9cc3ffff",
		16#4635# => X"90e60000",
		16#4636# => X"bc070039",
		16#4637# => X"0c0001ed",
		16#4638# => X"e4262000",
		16#4639# => X"13fffffa",
		16#463a# => X"15000000",
		16#463b# => X"84c10008",
		16#463c# => X"d4011828",
		16#463d# => X"9cc60001",
		16#463e# => X"9c600031",
		16#463f# => X"84e10020",
		16#4640# => X"d4013008",
		16#4641# => X"03fffe17",
		16#4642# => X"d8071800",
		16#4643# => X"e0ce3004",
		16#4644# => X"bd660000",
		16#4645# => X"13fffe1e",
		16#4646# => X"a87e0000",
		16#4647# => X"0400092f",
		16#4648# => X"a88e0000",
		16#4649# => X"03fffe1b",
		16#464a# => X"a87e0000",
		16#464b# => X"9d800020",
		16#464c# => X"e18c6802",
		16#464d# => X"bdac0004",
		16#464e# => X"1000022d",
		16#464f# => X"84c10034",
		16#4650# => X"9d8cfffc",
		16#4651# => X"e0846000",
		16#4652# => X"e0c66000",
		16#4653# => X"e1ce6000",
		16#4654# => X"d4013034",
		16#4655# => X"03fffe89",
		16#4656# => X"d4012024",
		16#4657# => X"84810008",
		16#4658# => X"e2002002",
		16#4659# => X"bc100000",
		16#465a# => X"13fffd77",
		16#465b# => X"9f400002",
		16#465c# => X"a5f0000f",
		16#465d# => X"18c00001",
		16#465e# => X"b9ef0003",
		16#465f# => X"86610010",
		16#4660# => X"a8c68b04",
		16#4661# => X"a99c0000",
		16#4662# => X"e1ef3000",
		16#4663# => X"a9b30000",
		16#4664# => X"e06c0004",
		16#4665# => X"e08d0004",
		16#4666# => X"84af0000",
		16#4667# => X"84cf0004",
		16#4668# => X"07ffe6a1",
		16#4669# => X"ba100084",
		16#466a# => X"d401602c",
		16#466b# => X"bc100000",
		16#466c# => X"13fffd65",
		16#466d# => X"aa4b0000",
		16#466e# => X"1a800001",
		16#466f# => X"a9d20000",
		16#4670# => X"aa948bcc",
		16#4671# => X"a9ac0000",
		16#4672# => X"a9720000",
		16#4673# => X"a4500001",
		16#4674# => X"a86e0000",
		16#4675# => X"a88d0000",
		16#4676# => X"bc020000",
		16#4677# => X"10000006",
		16#4678# => X"ba100081",
		16#4679# => X"84b40000",
		16#467a# => X"84d40004",
		16#467b# => X"07ffe68e",
		16#467c# => X"9f5a0001",
		16#467d# => X"a9cb0000",
		16#467e# => X"a9ac0000",
		16#467f# => X"bc300000",
		16#4680# => X"13fffff3",
		16#4681# => X"9e940008",
		16#4682# => X"aa4b0000",
		16#4683# => X"03fffd4e",
		16#4684# => X"d401602c",
		16#4685# => X"18c00001",
		16#4686# => X"9c84ffff",
		16#4687# => X"a8c68b04",
		16#4688# => X"b9840003",
		16#4689# => X"aaee0000",
		16#468a# => X"aada0000",
		16#468b# => X"e18c3000",
		16#468c# => X"d4012050",
		16#468d# => X"e0b60004",
		16#468e# => X"e0d70004",
		16#468f# => X"846c0000",
		16#4690# => X"848c0004",
		16#4691# => X"07ffe678",
		16#4692# => X"aa920000",
		16#4693# => X"8461002c",
		16#4694# => X"84e10020",
		16#4695# => X"aaa30000",
		16#4696# => X"9ce70001",
		16#4697# => X"e0740004",
		16#4698# => X"e0950004",
		16#4699# => X"d4013828",
		16#469a# => X"d4016060",
		16#469b# => X"07ffe9d9",
		16#469c# => X"d4015854",
		16#469d# => X"a86b0000",
		16#469e# => X"07ffe951",
		16#469f# => X"a9cb0000",
		16#46a0# => X"85e1002c",
		16#46a1# => X"e0ab0004",
		16#46a2# => X"e0cc0004",
		16#46a3# => X"aaaf0000",
		16#46a4# => X"e0740004",
		16#46a5# => X"e0950004",
		16#46a6# => X"07ffe641",
		16#46a7# => X"15000000",
		16#46a8# => X"9dae0030",
		16#46a9# => X"84610020",
		16#46aa# => X"8441004c",
		16#46ab# => X"d8036800",
		16#46ac# => X"aacb0000",
		16#46ad# => X"bc220001",
		16#46ae# => X"0c00002a",
		16#46af# => X"aa8c0000",
		16#46b0# => X"84c10020",
		16#46b1# => X"84e1004c",
		16#46b2# => X"87410028",
		16#46b3# => X"e2463800",
		16#46b4# => X"a9760000",
		16#46b5# => X"18400001",
		16#46b6# => X"a86b0000",
		16#46b7# => X"a8428a9c",
		16#46b8# => X"84a20000",
		16#46b9# => X"84c20004",
		16#46ba# => X"07ffe64f",
		16#46bb# => X"a88c0000",
		16#46bc# => X"aa0b0000",
		16#46bd# => X"a88c0000",
		16#46be# => X"a8700000",
		16#46bf# => X"07ffe9b5",
		16#46c0# => X"a9cc0000",
		16#46c1# => X"a86b0000",
		16#46c2# => X"07ffe92d",
		16#46c3# => X"aa8b0000",
		16#46c4# => X"a8500000",
		16#46c5# => X"a86e0000",
		16#46c6# => X"e0ab0004",
		16#46c7# => X"e0cc0004",
		16#46c8# => X"e0830004",
		16#46c9# => X"e0620004",
		16#46ca# => X"07ffe61d",
		16#46cb# => X"15000000",
		16#46cc# => X"9c740030",
		16#46cd# => X"d81a1800",
		16#46ce# => X"9f5a0001",
		16#46cf# => X"e43a9000",
		16#46d0# => X"13ffffe6",
		16#46d1# => X"18400001",
		16#46d2# => X"84610028",
		16#46d3# => X"84810050",
		16#46d4# => X"aacb0000",
		16#46d5# => X"e0632000",
		16#46d6# => X"aa8c0000",
		16#46d7# => X"d4011828",
		16#46d8# => X"85a10054",
		16#46d9# => X"84610060",
		16#46da# => X"19c00001",
		16#46db# => X"a9ed0000",
		16#46dc# => X"aa030000",
		16#46dd# => X"a9ce8ab4",
		16#46de# => X"e06f0004",
		16#46df# => X"e0900004",
		16#46e0# => X"84ae0000",
		16#46e1# => X"84ce0004",
		16#46e2# => X"07ffe5e6",
		16#46e3# => X"aa140000",
		16#46e4# => X"a9f60000",
		16#46e5# => X"e0ab0004",
		16#46e6# => X"e0cc0004",
		16#46e7# => X"e06f0004",
		16#46e8# => X"e0900004",
		16#46e9# => X"07ffe872",
		16#46ea# => X"15000000",
		16#46eb# => X"bd4b0000",
		16#46ec# => X"13fffc60",
		16#46ed# => X"84610028",
		16#46ee# => X"85810060",
		16#46ef# => X"84410054",
		16#46f0# => X"aa0c0000",
		16#46f1# => X"a9e20000",
		16#46f2# => X"846e0000",
		16#46f3# => X"848e0004",
		16#46f4# => X"e0af0004",
		16#46f5# => X"e0d00004",
		16#46f6# => X"07ffe5f1",
		16#46f7# => X"a9d60000",
		16#46f8# => X"a9f40000",
		16#46f9# => X"e0ab0004",
		16#46fa# => X"e0cc0004",
		16#46fb# => X"e06e0004",
		16#46fc# => X"e08f0004",
		16#46fd# => X"07ffe89a",
		16#46fe# => X"15000000",
		16#46ff# => X"bd8b0000",
		16#4700# => X"0ffffb81",
		16#4701# => X"84c10008",
		16#4702# => X"00000003",
		16#4703# => X"84810028",
		16#4704# => X"a8820000",
		16#4705# => X"9c44ffff",
		16#4706# => X"90620000",
		16#4707# => X"bc030030",
		16#4708# => X"13fffffc",
		16#4709# => X"15000000",
		16#470a# => X"d4012028",
		16#470b# => X"8481005c",
		16#470c# => X"03fffd5a",
		16#470d# => X"d4012008",
		16#470e# => X"9c800000",
		16#470f# => X"03fffb4f",
		16#4710# => X"d4012044",
		16#4711# => X"9cc00001",
		16#4712# => X"d4013044",
		16#4713# => X"84410018",
		16#4714# => X"bda20000",
		16#4715# => X"1000002c",
		16#4716# => X"aa220000",
		16#4717# => X"d4011038",
		16#4718# => X"03fffb4e",
		16#4719# => X"d401101c",
		16#471a# => X"9ce00000",
		16#471b# => X"03fffff8",
		16#471c# => X"d4013844",
		16#471d# => X"84610030",
		16#471e# => X"04000aad",
		16#471f# => X"a8820000",
		16#4720# => X"bd6b0000",
		16#4721# => X"13fffdd4",
		16#4722# => X"84c1001c",
		16#4723# => X"84e10008",
		16#4724# => X"a87e0000",
		16#4725# => X"84810030",
		16#4726# => X"9ce7ffff",
		16#4727# => X"9ca0000a",
		16#4728# => X"9cc00000",
		16#4729# => X"04000859",
		16#472a# => X"d4013808",
		16#472b# => X"84610038",
		16#472c# => X"84810044",
		16#472d# => X"d4015830",
		16#472e# => X"bc040000",
		16#472f# => X"13fffdc5",
		16#4730# => X"d401181c",
		16#4731# => X"a8920000",
		16#4732# => X"a87e0000",
		16#4733# => X"9ca0000a",
		16#4734# => X"0400084e",
		16#4735# => X"9cc00000",
		16#4736# => X"03fffdbe",
		16#4737# => X"aa4b0000",
		16#4738# => X"85820010",
		16#4739# => X"9d8c0004",
		16#473a# => X"b98c0002",
		16#473b# => X"e1826000",
		16#473c# => X"040008d6",
		16#473d# => X"846c0000",
		16#473e# => X"9da00020",
		16#473f# => X"03fffd92",
		16#4740# => X"e1ad5802",
		16#4741# => X"9c600001",
		16#4742# => X"d4011838",
		16#4743# => X"d401181c",
		16#4744# => X"03fffc50",
		16#4745# => X"d4011818",
		16#4746# => X"bcb1000e",
		16#4747# => X"10000003",
		16#4748# => X"9d800001",
		16#4749# => X"9d800000",
		16#474a# => X"e1ce6003",
		16#474b# => X"03fffc49",
		16#474c# => X"d401881c",
		16#474d# => X"84e10010",
		16#474e# => X"e4278000",
		16#474f# => X"13fffd7f",
		16#4750# => X"84610048",
		16#4751# => X"1860000f",
		16#4752# => X"a863ffff",
		16#4753# => X"e19c1803",
		16#4754# => X"bc2c0000",
		16#4755# => X"13fffd78",
		16#4756# => X"aa070000",
		16#4757# => X"18807ff0",
		16#4758# => X"e39c2003",
		16#4759# => X"bc1c0000",
		16#475a# => X"13fffd74",
		16#475b# => X"84610048",
		16#475c# => X"84c10034",
		16#475d# => X"84e10024",
		16#475e# => X"9cc60001",
		16#475f# => X"9ce70001",
		16#4760# => X"d4013034",
		16#4761# => X"d4013824",
		16#4762# => X"03fffd6b",
		16#4763# => X"9e000001",
		16#4764# => X"10000006",
		16#4765# => X"a8920000",
		16#4766# => X"a87e0000",
		16#4767# => X"04000a05",
		16#4768# => X"a8ae0000",
		16#4769# => X"aa4b0000",
		16#476a# => X"bc100000",
		16#476b# => X"0c0000bd",
		16#476c# => X"aa920000",
		16#476d# => X"9f400001",
		16#476e# => X"84c10010",
		16#476f# => X"84810020",
		16#4770# => X"e386d003",
		16#4771# => X"d4012028",
		16#4772# => X"d401e018",
		16#4773# => X"a9d20000",
		16#4774# => X"ab9a0000",
		16#4775# => X"87010030",
		16#4776# => X"ab440000",
		16#4777# => X"a8780000",
		16#4778# => X"a8820000",
		16#4779# => X"07fff945",
		16#477a# => X"9ec00001",
		16#477b# => X"a8780000",
		16#477c# => X"a88e0000",
		16#477d# => X"9d6b0030",
		16#477e# => X"04000a4d",
		16#477f# => X"d4015810",
		16#4780# => X"a87e0000",
		16#4781# => X"a8820000",
		16#4782# => X"a8b40000",
		16#4783# => X"04000a63",
		16#4784# => X"aa0b0000",
		16#4785# => X"846b000c",
		16#4786# => X"bc230000",
		16#4787# => X"0c000035",
		16#4788# => X"aa4b0000",
		16#4789# => X"a87e0000",
		16#478a# => X"040007ec",
		16#478b# => X"a8920000",
		16#478c# => X"84e10000",
		16#478d# => X"e0763804",
		16#478e# => X"bc230000",
		16#478f# => X"10000006",
		16#4790# => X"bd900000",
		16#4791# => X"84610018",
		16#4792# => X"bc230000",
		16#4793# => X"0c0000c4",
		16#4794# => X"bd900000",
		16#4795# => X"10000067",
		16#4796# => X"84c10000",
		16#4797# => X"e2103004",
		16#4798# => X"bc300000",
		16#4799# => X"10000006",
		16#479a# => X"bdb60000",
		16#479b# => X"84e10018",
		16#479c# => X"bc270000",
		16#479d# => X"0c00005f",
		16#479e# => X"bdb60000",
		16#479f# => X"0c0000a3",
		16#47a0# => X"84610010",
		16#47a1# => X"d81a1800",
		16#47a2# => X"8481001c",
		16#47a3# => X"e41c2000",
		16#47a4# => X"10000099",
		16#47a5# => X"9f5a0001",
		16#47a6# => X"a8980000",
		16#47a7# => X"a87e0000",
		16#47a8# => X"9ca0000a",
		16#47a9# => X"040007d9",
		16#47aa# => X"9cc00000",
		16#47ab# => X"e42ea000",
		16#47ac# => X"0c000015",
		16#47ad# => X"ab0b0000",
		16#47ae# => X"a88e0000",
		16#47af# => X"9ca0000a",
		16#47b0# => X"9cc00000",
		16#47b1# => X"a87e0000",
		16#47b2# => X"040007d0",
		16#47b3# => X"9f9c0001",
		16#47b4# => X"a8940000",
		16#47b5# => X"a87e0000",
		16#47b6# => X"9ca0000a",
		16#47b7# => X"9cc00000",
		16#47b8# => X"040007ca",
		16#47b9# => X"a9cb0000",
		16#47ba# => X"03ffffbd",
		16#47bb# => X"aa8b0000",
		16#47bc# => X"a8780000",
		16#47bd# => X"04000a0e",
		16#47be# => X"a88b0000",
		16#47bf# => X"03ffffca",
		16#47c0# => X"aacb0000",
		16#47c1# => X"a88e0000",
		16#47c2# => X"a87e0000",
		16#47c3# => X"9ca0000a",
		16#47c4# => X"9cc00000",
		16#47c5# => X"040007bd",
		16#47c6# => X"9f9c0001",
		16#47c7# => X"a9cb0000",
		16#47c8# => X"03ffffaf",
		16#47c9# => X"aa8b0000",
		16#47ca# => X"03fffc9c",
		16#47cb# => X"d401b028",
		16#47cc# => X"a87e0000",
		16#47cd# => X"84810030",
		16#47ce# => X"04000946",
		16#47cf# => X"84a10040",
		16#47d0# => X"03fffced",
		16#47d1# => X"d4015830",
		16#47d2# => X"84610048",
		16#47d3# => X"e1901002",
		16#47d4# => X"9e000000",
		16#47d5# => X"e0636000",
		16#47d6# => X"e0426000",
		16#47d7# => X"d4011848",
		16#47d8# => X"03fffcaa",
		16#47d9# => X"d4011040",
		16#47da# => X"84810030",
		16#47db# => X"04000939",
		16#47dc# => X"a8b00000",
		16#47dd# => X"03fffce0",
		16#47de# => X"d4015830",
		16#47df# => X"9c400000",
		16#47e0# => X"03fffc72",
		16#47e1# => X"aa420000",
		16#47e2# => X"84810058",
		16#47e3# => X"bc040000",
		16#47e4# => X"10000054",
		16#47e5# => X"9c400036",
		16#47e6# => X"9dad0433",
		16#47e7# => X"86010040",
		16#47e8# => X"03fffca0",
		16#47e9# => X"85c10034",
		16#47ea# => X"9cc60001",
		16#47eb# => X"d4011828",
		16#47ec# => X"b8c60018",
		16#47ed# => X"8461005c",
		16#47ee# => X"d4012020",
		16#47ef# => X"b8c60098",
		16#47f0# => X"d4011808",
		16#47f1# => X"03fffc75",
		16#47f2# => X"d8023000",
		16#47f3# => X"84810020",
		16#47f4# => X"03fffb5b",
		16#47f5# => X"87c10060",
		16#47f6# => X"87c10060",
		16#47f7# => X"03fffa89",
		16#47f8# => X"87810064",
		16#47f9# => X"9da00000",
		16#47fa# => X"03fffc8e",
		16#47fb# => X"e1c62002",
		16#47fc# => X"d401c030",
		16#47fd# => X"d401d028",
		16#47fe# => X"bdb60000",
		16#47ff# => X"1000000f",
		16#4800# => X"86010010",
		16#4801# => X"9ca00001",
		16#4802# => X"a87e0000",
		16#4803# => X"04000969",
		16#4804# => X"a8980000",
		16#4805# => X"a8820000",
		16#4806# => X"a86b0000",
		16#4807# => X"040009c4",
		16#4808# => X"d4015830",
		16#4809# => X"bd4b0000",
		16#480a# => X"0c00005d",
		16#480b# => X"bc100039",
		16#480c# => X"10000042",
		16#480d# => X"9e100001",
		16#480e# => X"84610028",
		16#480f# => X"aa540000",
		16#4810# => X"d8038000",
		16#4811# => X"9c630001",
		16#4812# => X"03fffc46",
		16#4813# => X"d4011828",
		16#4814# => X"10000009",
		16#4815# => X"84a10028",
		16#4816# => X"a6100001",
		16#4817# => X"bc300000",
		16#4818# => X"13fffe19",
		16#4819# => X"84610028",
		16#481a# => X"00000004",
		16#481b# => X"9c65ffff",
		16#481c# => X"a8a30000",
		16#481d# => X"9c65ffff",
		16#481e# => X"90830000",
		16#481f# => X"bc040030",
		16#4820# => X"13fffffc",
		16#4821# => X"15000000",
		16#4822# => X"03fffc36",
		16#4823# => X"d4012828",
		16#4824# => X"9ce70001",
		16#4825# => X"d4011828",
		16#4826# => X"03fffc32",
		16#4827# => X"d8063800",
		16#4828# => X"a87e0000",
		16#4829# => X"04000720",
		16#482a# => X"84920004",
		16#482b# => X"84f20010",
		16#482c# => X"9c6b000c",
		16#482d# => X"9ce70002",
		16#482e# => X"9c92000c",
		16#482f# => X"b8a70002",
		16#4830# => X"04000626",
		16#4831# => X"a9cb0000",
		16#4832# => X"a87e0000",
		16#4833# => X"a88e0000",
		16#4834# => X"04000938",
		16#4835# => X"9ca00001",
		16#4836# => X"03ffff37",
		16#4837# => X"aa8b0000",
		16#4838# => X"85a1006c",
		16#4839# => X"86010040",
		16#483a# => X"e1a26802",
		16#483b# => X"03fffc4d",
		16#483c# => X"85c10034",
		16#483d# => X"86010010",
		16#483e# => X"d401c030",
		16#483f# => X"d401d028",
		16#4840# => X"03fffde5",
		16#4841# => X"aa540000",
		16#4842# => X"86010010",
		16#4843# => X"d401c030",
		16#4844# => X"bc300039",
		16#4845# => X"0c000009",
		16#4846# => X"d401d028",
		16#4847# => X"84e10028",
		16#4848# => X"9e100001",
		16#4849# => X"aa540000",
		16#484a# => X"d8078000",
		16#484b# => X"9ce70001",
		16#484c# => X"03fffc0c",
		16#484d# => X"d4013828",
		16#484e# => X"84810028",
		16#484f# => X"9cc00039",
		16#4850# => X"aa540000",
		16#4851# => X"d8043000",
		16#4852# => X"9c840001",
		16#4853# => X"d4012028",
		16#4854# => X"a8640000",
		16#4855# => X"03fffddf",
		16#4856# => X"84810020",
		16#4857# => X"d401c030",
		16#4858# => X"d401d028",
		16#4859# => X"ab100000",
		16#485a# => X"86010010",
		16#485b# => X"bc100039",
		16#485c# => X"13fffff2",
		16#485d# => X"bdb80000",
		16#485e# => X"10000003",
		16#485f# => X"15000000",
		16#4860# => X"9e100001",
		16#4861# => X"84810028",
		16#4862# => X"aa540000",
		16#4863# => X"d8048000",
		16#4864# => X"9c840001",
		16#4865# => X"03fffbf3",
		16#4866# => X"d4012028",
		16#4867# => X"bc2b0000",
		16#4868# => X"13ffffa7",
		16#4869# => X"84610028",
		16#486a# => X"a4700001",
		16#486b# => X"bc030000",
		16#486c# => X"13ffffa3",
		16#486d# => X"84610028",
		16#486e# => X"03ffff9e",
		16#486f# => X"bc100039",
		16#4870# => X"8481005c",
		16#4871# => X"03fffbf5",
		16#4872# => X"d4012008",
		16#4873# => X"8461001c",
		16#4874# => X"bca3000e",
		16#4875# => X"10000003",
		16#4876# => X"9c400001",
		16#4877# => X"9c400000",
		16#4878# => X"e1ce1003",
		16#4879# => X"03fffb1d",
		16#487a# => X"9c400000",
		16#487b# => X"bc0c0004",
		16#487c# => X"13fffc63",
		16#487d# => X"84810034",
		16#487e# => X"03fffc59",
		16#487f# => X"9d8c001c",
		16#4880# => X"d7e117ec",
		16#4881# => X"d7e197f8",
		16#4882# => X"d7e14ffc",
		16#4883# => X"d7e177f0",
		16#4884# => X"d7e187f4",
		16#4885# => X"aa430000",
		16#4886# => X"9c21ffec",
		16#4887# => X"bc030000",
		16#4888# => X"10000006",
		16#4889# => X"a8440000",
		16#488a# => X"84830038",
		16#488b# => X"bc240000",
		16#488c# => X"0c00007b",
		16#488d# => X"15000000",
		16#488e# => X"9962000c",
		16#488f# => X"bc0b0000",
		16#4890# => X"10000048",
		16#4891# => X"a88b0000",
		16#4892# => X"a46b0008",
		16#4893# => X"bc230000",
		16#4894# => X"1000004b",
		16#4895# => X"15000000",
		16#4896# => X"a88b0800",
		16#4897# => X"84a20004",
		16#4898# => X"bd450000",
		16#4899# => X"0c000086",
		16#489a# => X"dc02200c",
		16#489b# => X"84e20028",
		16#489c# => X"bc070000",
		16#489d# => X"1000003b",
		16#489e# => X"a9670000",
		16#489f# => X"a464ffff",
		16#48a0# => X"9c800000",
		16#48a1# => X"85d20000",
		16#48a2# => X"a4a31000",
		16#48a3# => X"e4052000",
		16#48a4# => X"10000069",
		16#48a5# => X"d4122000",
		16#48a6# => X"84a20050",
		16#48a7# => X"a4630004",
		16#48a8# => X"bc030000",
		16#48a9# => X"1000000a",
		16#48aa# => X"a8720000",
		16#48ab# => X"84820004",
		16#48ac# => X"84620030",
		16#48ad# => X"bc030000",
		16#48ae# => X"10000004",
		16#48af# => X"e0a52002",
		16#48b0# => X"8462003c",
		16#48b1# => X"e0a51802",
		16#48b2# => X"a8720000",
		16#48b3# => X"8482001c",
		16#48b4# => X"48003800",
		16#48b5# => X"9cc00000",
		16#48b6# => X"bc2bffff",
		16#48b7# => X"0c00006e",
		16#48b8# => X"15000000",
		16#48b9# => X"9462000c",
		16#48ba# => X"9ca0f7ff",
		16#48bb# => X"84820010",
		16#48bc# => X"e0632803",
		16#48bd# => X"9ca00000",
		16#48be# => X"b8630010",
		16#48bf# => X"d4022000",
		16#48c0# => X"d4022804",
		16#48c1# => X"b8630090",
		16#48c2# => X"a4831000",
		16#48c3# => X"e4042800",
		16#48c4# => X"10000006",
		16#48c5# => X"dc02180c",
		16#48c6# => X"bc2bffff",
		16#48c7# => X"0c00006a",
		16#48c8# => X"15000000",
		16#48c9# => X"d4025850",
		16#48ca# => X"84820030",
		16#48cb# => X"d4127000",
		16#48cc# => X"bc040000",
		16#48cd# => X"1000000b",
		16#48ce# => X"a9640000",
		16#48cf# => X"9c620040",
		16#48d0# => X"e4041800",
		16#48d1# => X"10000005",
		16#48d2# => X"9c600000",
		16#48d3# => X"040001dc",
		16#48d4# => X"a8720000",
		16#48d5# => X"9c600000",
		16#48d6# => X"d4021830",
		16#48d7# => X"a9630000",
		16#48d8# => X"9c210014",
		16#48d9# => X"8521fffc",
		16#48da# => X"8441ffec",
		16#48db# => X"85c1fff0",
		16#48dc# => X"8601fff4",
		16#48dd# => X"44004800",
		16#48de# => X"8641fff8",
		16#48df# => X"85c20010",
		16#48e0# => X"bc0e0000",
		16#48e1# => X"13fffff7",
		16#48e2# => X"a96e0000",
		16#48e3# => X"86020000",
		16#48e4# => X"a4840003",
		16#48e5# => X"9c600000",
		16#48e6# => X"d4027000",
		16#48e7# => X"e4241800",
		16#48e8# => X"0c000023",
		16#48e9# => X"e2107002",
		16#48ea# => X"9d600000",
		16#48eb# => X"e5b05800",
		16#48ec# => X"0c000007",
		16#48ed# => X"d4021808",
		16#48ee# => X"03ffffeb",
		16#48ef# => X"9c210014",
		16#48f0# => X"bdb00000",
		16#48f1# => X"10000026",
		16#48f2# => X"e1ce5800",
		16#48f3# => X"a8d00000",
		16#48f4# => X"a8ae0000",
		16#48f5# => X"85620024",
		16#48f6# => X"a8720000",
		16#48f7# => X"48005800",
		16#48f8# => X"8482001c",
		16#48f9# => X"bd4b0000",
		16#48fa# => X"13fffff6",
		16#48fb# => X"e2105802",
		16#48fc# => X"9462000c",
		16#48fd# => X"a8630040",
		16#48fe# => X"9d60ffff",
		16#48ff# => X"dc02180c",
		16#4900# => X"9c210014",
		16#4901# => X"8521fffc",
		16#4902# => X"8441ffec",
		16#4903# => X"85c1fff0",
		16#4904# => X"8601fff4",
		16#4905# => X"44004800",
		16#4906# => X"8641fff8",
		16#4907# => X"04000087",
		16#4908# => X"15000000",
		16#4909# => X"03ffff86",
		16#490a# => X"9962000c",
		16#490b# => X"03ffffdf",
		16#490c# => X"84620014",
		16#490d# => X"a8720000",
		16#490e# => X"8482001c",
		16#490f# => X"48003800",
		16#4910# => X"9cc00001",
		16#4911# => X"bc2bffff",
		16#4912# => X"0c000025",
		16#4913# => X"a8ab0000",
		16#4914# => X"9462000c",
		16#4915# => X"03ffff92",
		16#4916# => X"84e20028",
		16#4917# => X"9c210014",
		16#4918# => X"9d600000",
		16#4919# => X"8521fffc",
		16#491a# => X"8441ffec",
		16#491b# => X"85c1fff0",
		16#491c# => X"8601fff4",
		16#491d# => X"44004800",
		16#491e# => X"8641fff8",
		16#491f# => X"84a2003c",
		16#4920# => X"bda50000",
		16#4921# => X"0fffff7a",
		16#4922# => X"a9630000",
		16#4923# => X"03ffffb6",
		16#4924# => X"9c210014",
		16#4925# => X"84720000",
		16#4926# => X"bc030000",
		16#4927# => X"13ffff92",
		16#4928# => X"bc03001d",
		16#4929# => X"13ffff90",
		16#492a# => X"bc230016",
		16#492b# => X"0fffff8e",
		16#492c# => X"15000000",
		16#492d# => X"9462000c",
		16#492e# => X"a8630040",
		16#492f# => X"03ffffa9",
		16#4930# => X"dc02180c",
		16#4931# => X"84720000",
		16#4932# => X"e4232800",
		16#4933# => X"13ffff97",
		16#4934# => X"15000000",
		16#4935# => X"03ffff95",
		16#4936# => X"d4025850",
		16#4937# => X"84720000",
		16#4938# => X"bc230000",
		16#4939# => X"0fffffdb",
		16#493a# => X"ac830016",
		16#493b# => X"e0c02002",
		16#493c# => X"e0862004",
		16#493d# => X"bd640000",
		16#493e# => X"10000007",
		16#493f# => X"ac63001d",
		16#4940# => X"e0801802",
		16#4941# => X"e0641804",
		16#4942# => X"bd830000",
		16#4943# => X"10000005",
		16#4944# => X"15000000",
		16#4945# => X"d4127000",
		16#4946# => X"03ffff92",
		16#4947# => X"9d600000",
		16#4948# => X"9462000c",
		16#4949# => X"a8630040",
		16#494a# => X"03ffff8e",
		16#494b# => X"dc02180c",
		16#494c# => X"d7e14ffc",
		16#494d# => X"bc230000",
		16#494e# => X"0c00000a",
		16#494f# => X"9c21fffc",
		16#4950# => X"a8830000",
		16#4951# => X"18600001",
		16#4952# => X"a863ade4",
		16#4953# => X"84630000",
		16#4954# => X"9c210004",
		16#4955# => X"8521fffc",
		16#4956# => X"03ffff2a",
		16#4957# => X"15000000",
		16#4958# => X"18600001",
		16#4959# => X"18800001",
		16#495a# => X"a8638890",
		16#495b# => X"9c210004",
		16#495c# => X"a8842200",
		16#495d# => X"8521fffc",
		16#495e# => X"000003c0",
		16#495f# => X"84630000",
		16#4960# => X"44004800",
		16#4961# => X"9d600000",
		16#4962# => X"44004800",
		16#4963# => X"9d600000",
		16#4964# => X"d7e14ffc",
		16#4965# => X"9c21fffc",
		16#4966# => X"18800001",
		16#4967# => X"9c210004",
		16#4968# => X"8521fffc",
		16#4969# => X"00000383",
		16#496a# => X"a8847064",
		16#496b# => X"d7e177f4",
		16#496c# => X"9dc00068",
		16#496d# => X"d7e117f0",
		16#496e# => X"e1c47306",
		16#496f# => X"d7e187f8",
		16#4970# => X"d7e14ffc",
		16#4971# => X"aa040000",
		16#4972# => X"9c21fff0",
		16#4973# => X"07ffe817",
		16#4974# => X"9c8e000c",
		16#4975# => X"bc0b0000",
		16#4976# => X"10000009",
		16#4977# => X"a84b0000",
		16#4978# => X"9c6b000c",
		16#4979# => X"9c800000",
		16#497a# => X"d40b8004",
		16#497b# => X"d40b2000",
		16#497c# => X"d40b1808",
		16#497d# => X"0400057c",
		16#497e# => X"a8ae0000",
		16#497f# => X"9c210010",
		16#4980# => X"a9620000",
		16#4981# => X"8521fffc",
		16#4982# => X"8441fff0",
		16#4983# => X"85c1fff4",
		16#4984# => X"44004800",
		16#4985# => X"8601fff8",
		16#4986# => X"d7e14ffc",
		16#4987# => X"18600001",
		16#4988# => X"9c21fffc",
		16#4989# => X"a8638890",
		16#498a# => X"9c210004",
		16#498b# => X"8521fffc",
		16#498c# => X"03ffffd8",
		16#498d# => X"84630000",
		16#498e# => X"d7e117d8",
		16#498f# => X"d7e197e4",
		16#4990# => X"d7e14ffc",
		16#4991# => X"d7e177dc",
		16#4992# => X"d7e187e0",
		16#4993# => X"d7e1a7e8",
		16#4994# => X"d7e1b7ec",
		16#4995# => X"d7e1c7f0",
		16#4996# => X"d7e1d7f4",
		16#4997# => X"d7e1e7f8",
		16#4998# => X"84430038",
		16#4999# => X"9c21ffd8",
		16#499a# => X"bc220000",
		16#499b# => X"10000051",
		16#499c# => X"aa430000",
		16#499d# => X"18800001",
		16#499e# => X"9f800001",
		16#499f# => X"a8842590",
		16#49a0# => X"9c6302ec",
		16#49a1# => X"d412203c",
		16#49a2# => X"9c800003",
		16#49a3# => X"85d20004",
		16#49a4# => X"9cc00004",
		16#49a5# => X"d41222e4",
		16#49a6# => X"d4121ae8",
		16#49a7# => X"d412e038",
		16#49a8# => X"d41212e0",
		16#49a9# => X"9c6e005c",
		16#49aa# => X"dc0e300c",
		16#49ab# => X"a8820000",
		16#49ac# => X"9ca00008",
		16#49ad# => X"d40e1000",
		16#49ae# => X"d40e1004",
		16#49af# => X"d40e1008",
		16#49b0# => X"d40e1064",
		16#49b1# => X"dc0e100e",
		16#49b2# => X"d40e1010",
		16#49b3# => X"d40e1014",
		16#49b4# => X"d40e1018",
		16#49b5# => X"1b400001",
		16#49b6# => X"1b000001",
		16#49b7# => X"1ac00001",
		16#49b8# => X"04000541",
		16#49b9# => X"1a800001",
		16#49ba# => X"ab5a59dc",
		16#49bb# => X"86120008",
		16#49bc# => X"ab185a40",
		16#49bd# => X"aad65ac4",
		16#49be# => X"aa945b24",
		16#49bf# => X"9cc00009",
		16#49c0# => X"9c70005c",
		16#49c1# => X"a8820000",
		16#49c2# => X"9ca00008",
		16#49c3# => X"d40e701c",
		16#49c4# => X"d40ed020",
		16#49c5# => X"d40ec024",
		16#49c6# => X"d40eb028",
		16#49c7# => X"d40ea02c",
		16#49c8# => X"dc10300c",
		16#49c9# => X"d4101000",
		16#49ca# => X"d4101004",
		16#49cb# => X"d4101008",
		16#49cc# => X"d4101064",
		16#49cd# => X"dc10e00e",
		16#49ce# => X"d4101010",
		16#49cf# => X"d4101014",
		16#49d0# => X"04000529",
		16#49d1# => X"d4101018",
		16#49d2# => X"9c600012",
		16#49d3# => X"85d2000c",
		16#49d4# => X"9cc00002",
		16#49d5# => X"dc0e180c",
		16#49d6# => X"d410801c",
		16#49d7# => X"d410d020",
		16#49d8# => X"d410c024",
		16#49d9# => X"d410b028",
		16#49da# => X"d410a02c",
		16#49db# => X"d40e1000",
		16#49dc# => X"d40e1004",
		16#49dd# => X"d40e1008",
		16#49de# => X"d40e1064",
		16#49df# => X"dc0e300e",
		16#49e0# => X"d40e1010",
		16#49e1# => X"d40e1014",
		16#49e2# => X"d40e1018",
		16#49e3# => X"9c6e005c",
		16#49e4# => X"a8820000",
		16#49e5# => X"04000514",
		16#49e6# => X"9ca00008",
		16#49e7# => X"d40e701c",
		16#49e8# => X"d40ed020",
		16#49e9# => X"d40ec024",
		16#49ea# => X"d40eb028",
		16#49eb# => X"d40ea02c",
		16#49ec# => X"9c210028",
		16#49ed# => X"8521fffc",
		16#49ee# => X"8441ffd8",
		16#49ef# => X"85c1ffdc",
		16#49f0# => X"8601ffe0",
		16#49f1# => X"8641ffe4",
		16#49f2# => X"8681ffe8",
		16#49f3# => X"86c1ffec",
		16#49f4# => X"8701fff0",
		16#49f5# => X"8741fff4",
		16#49f6# => X"44004800",
		16#49f7# => X"8781fff8",
		16#49f8# => X"d7e117f0",
		16#49f9# => X"18400001",
		16#49fa# => X"d7e177f4",
		16#49fb# => X"a8428890",
		16#49fc# => X"d7e187f8",
		16#49fd# => X"85c20000",
		16#49fe# => X"d7e14ffc",
		16#49ff# => X"844e0038",
		16#4a00# => X"9c21fff0",
		16#4a01# => X"bc220000",
		16#4a02# => X"0c000033",
		16#4a03# => X"aa030000",
		16#4a04# => X"9dce02e0",
		16#4a05# => X"848e0004",
		16#4a06# => X"9c84ffff",
		16#4a07# => X"bd840000",
		16#4a08# => X"0c000007",
		16#4a09# => X"844e0008",
		16#4a0a# => X"00000026",
		16#4a0b# => X"856e0000",
		16#4a0c# => X"bd640000",
		16#4a0d# => X"0c000022",
		16#4a0e# => X"9c420068",
		16#4a0f# => X"98a2000c",
		16#4a10# => X"bc050000",
		16#4a11# => X"0ffffffb",
		16#4a12# => X"9c84ffff",
		16#4a13# => X"9c60ffff",
		16#4a14# => X"9c800000",
		16#4a15# => X"dc02180e",
		16#4a16# => X"9c600001",
		16#4a17# => X"9ca00008",
		16#4a18# => X"dc02180c",
		16#4a19# => X"9c600000",
		16#4a1a# => X"d4021864",
		16#4a1b# => X"d4021800",
		16#4a1c# => X"d4021808",
		16#4a1d# => X"d4021804",
		16#4a1e# => X"d4021810",
		16#4a1f# => X"d4021814",
		16#4a20# => X"d4021818",
		16#4a21# => X"040004d8",
		16#4a22# => X"9c62005c",
		16#4a23# => X"9c600000",
		16#4a24# => X"d4021830",
		16#4a25# => X"d4021834",
		16#4a26# => X"d4021844",
		16#4a27# => X"d4021848",
		16#4a28# => X"9c210010",
		16#4a29# => X"a9620000",
		16#4a2a# => X"8521fffc",
		16#4a2b# => X"8441fff0",
		16#4a2c# => X"85c1fff4",
		16#4a2d# => X"44004800",
		16#4a2e# => X"8601fff8",
		16#4a2f# => X"856e0000",
		16#4a30# => X"bc2b0000",
		16#4a31# => X"0c000008",
		16#4a32# => X"15000000",
		16#4a33# => X"03ffffd2",
		16#4a34# => X"a9cb0000",
		16#4a35# => X"07ffff59",
		16#4a36# => X"a86e0000",
		16#4a37# => X"03ffffce",
		16#4a38# => X"9dce02e0",
		16#4a39# => X"a8700000",
		16#4a3a# => X"07ffff31",
		16#4a3b# => X"9c800004",
		16#4a3c# => X"bc0b0000",
		16#4a3d# => X"0ffffff6",
		16#4a3e# => X"d40e5800",
		16#4a3f# => X"9c60000c",
		16#4a40# => X"a84b0000",
		16#4a41# => X"03ffffe7",
		16#4a42# => X"d4101800",
		16#4a43# => X"44004800",
		16#4a44# => X"15000000",
		16#4a45# => X"44004800",
		16#4a46# => X"15000000",
		16#4a47# => X"44004800",
		16#4a48# => X"15000000",
		16#4a49# => X"44004800",
		16#4a4a# => X"15000000",
		16#4a4b# => X"18600001",
		16#4a4c# => X"d7e14ffc",
		16#4a4d# => X"a863ade4",
		16#4a4e# => X"9c21fffc",
		16#4a4f# => X"18800001",
		16#4a50# => X"84630000",
		16#4a51# => X"9c210004",
		16#4a52# => X"8521fffc",
		16#4a53# => X"00000299",
		16#4a54# => X"a8842580",
		16#4a55# => X"18600001",
		16#4a56# => X"d7e14ffc",
		16#4a57# => X"a863ade4",
		16#4a58# => X"9c21fffc",
		16#4a59# => X"18800001",
		16#4a5a# => X"84630000",
		16#4a5b# => X"9c210004",
		16#4a5c# => X"8521fffc",
		16#4a5d# => X"0000028f",
		16#4a5e# => X"a8842588",
		16#4a5f# => X"d7e117ec",
		16#4a60# => X"18400001",
		16#4a61# => X"d7e177f0",
		16#4a62# => X"d7e187f4",
		16#4a63# => X"d7e197f8",
		16#4a64# => X"d7e14ffc",
		16#4a65# => X"9c21ffec",
		16#4a66# => X"a842b20c",
		16#4a67# => X"aa440000",
		16#4a68# => X"07ffe972",
		16#4a69# => X"a9c30000",
		16#4a6a# => X"84620008",
		16#4a6b# => X"86030004",
		16#4a6c# => X"9c60fffc",
		16#4a6d# => X"e2101803",
		16#4a6e# => X"9c700fef",
		16#4a6f# => X"e2439002",
		16#4a70# => X"9c60f000",
		16#4a71# => X"e2521803",
		16#4a72# => X"e2521800",
		16#4a73# => X"bd520fff",
		16#4a74# => X"0c000009",
		16#4a75# => X"a86e0000",
		16#4a76# => X"07ffebf5",
		16#4a77# => X"9c800000",
		16#4a78# => X"84620008",
		16#4a79# => X"e0638000",
		16#4a7a# => X"e40b1800",
		16#4a7b# => X"1000000c",
		16#4a7c# => X"a86e0000",
		16#4a7d# => X"07ffe95f",
		16#4a7e# => X"a86e0000",
		16#4a7f# => X"9c210014",
		16#4a80# => X"9d600000",
		16#4a81# => X"8521fffc",
		16#4a82# => X"8441ffec",
		16#4a83# => X"85c1fff0",
		16#4a84# => X"8601fff4",
		16#4a85# => X"44004800",
		16#4a86# => X"8641fff8",
		16#4a87# => X"07ffebe4",
		16#4a88# => X"e0809002",
		16#4a89# => X"bc2bffff",
		16#4a8a# => X"0c000014",
		16#4a8b# => X"18800001",
		16#4a8c# => X"e2109002",
		16#4a8d# => X"a884c4c8",
		16#4a8e# => X"84420008",
		16#4a8f# => X"84640000",
		16#4a90# => X"aa100001",
		16#4a91# => X"e2439002",
		16#4a92# => X"d4028004",
		16#4a93# => X"a86e0000",
		16#4a94# => X"07ffe948",
		16#4a95# => X"d4049000",
		16#4a96# => X"9c210014",
		16#4a97# => X"9d600001",
		16#4a98# => X"8521fffc",
		16#4a99# => X"8441ffec",
		16#4a9a# => X"85c1fff0",
		16#4a9b# => X"8601fff4",
		16#4a9c# => X"44004800",
		16#4a9d# => X"8641fff8",
		16#4a9e# => X"a86e0000",
		16#4a9f# => X"07ffebcc",
		16#4aa0# => X"9c800000",
		16#4aa1# => X"84420008",
		16#4aa2# => X"e06b1002",
		16#4aa3# => X"bda3000f",
		16#4aa4# => X"13ffffd9",
		16#4aa5# => X"18800001",
		16#4aa6# => X"a8630001",
		16#4aa7# => X"a884b618",
		16#4aa8# => X"d4021804",
		16#4aa9# => X"84840000",
		16#4aaa# => X"18400001",
		16#4aab# => X"e16b2002",
		16#4aac# => X"a842c4c8",
		16#4aad# => X"03ffffd0",
		16#4aae# => X"d4025800",
		16#4aaf# => X"d7e117f4",
		16#4ab0# => X"d7e177f8",
		16#4ab1# => X"d7e14ffc",
		16#4ab2# => X"a9c40000",
		16#4ab3# => X"9c21fff4",
		16#4ab4# => X"bc040000",
		16#4ab5# => X"10000062",
		16#4ab6# => X"a8430000",
		16#4ab7# => X"07ffe923",
		16#4ab8# => X"15000000",
		16#4ab9# => X"9c8efff8",
		16#4aba# => X"9c60fffe",
		16#4abb# => X"18e00001",
		16#4abc# => X"85040004",
		16#4abd# => X"a8e7b20c",
		16#4abe# => X"e0a81803",
		16#4abf# => X"85670008",
		16#4ac0# => X"e0c42800",
		16#4ac1# => X"84660004",
		16#4ac2# => X"e42b3000",
		16#4ac3# => X"9d60fffc",
		16#4ac4# => X"0c00007c",
		16#4ac5# => X"e0635803",
		16#4ac6# => X"a5080001",
		16#4ac7# => X"9d600000",
		16#4ac8# => X"e4285800",
		16#4ac9# => X"1000000f",
		16#4aca# => X"d4061804",
		16#4acb# => X"85840000",
		16#4acc# => X"19a00001",
		16#4acd# => X"e0846002",
		16#4ace# => X"e0a56000",
		16#4acf# => X"a9adb214",
		16#4ad0# => X"85840008",
		16#4ad1# => X"e40c6800",
		16#4ad2# => X"10000006",
		16#4ad3# => X"9d600001",
		16#4ad4# => X"85a4000c",
		16#4ad5# => X"a9680000",
		16#4ad6# => X"d40c680c",
		16#4ad7# => X"d40d6008",
		16#4ad8# => X"e1061800",
		16#4ad9# => X"85080004",
		16#4ada# => X"a5080001",
		16#4adb# => X"bc280000",
		16#4adc# => X"10000008",
		16#4add# => X"bc2b0000",
		16#4ade# => X"0c00003e",
		16#4adf# => X"e0a51800",
		16#4ae0# => X"84660008",
		16#4ae1# => X"84c6000c",
		16#4ae2# => X"d403300c",
		16#4ae3# => X"d4061808",
		16#4ae4# => X"a8c50001",
		16#4ae5# => X"e0642800",
		16#4ae6# => X"d4043004",
		16#4ae7# => X"bc2b0000",
		16#4ae8# => X"10000029",
		16#4ae9# => X"d4032800",
		16#4aea# => X"bc4501ff",
		16#4aeb# => X"0c000040",
		16#4aec# => X"9cc00001",
		16#4aed# => X"b8650049",
		16#4aee# => X"bc430004",
		16#4aef# => X"1000006b",
		16#4af0# => X"bc430014",
		16#4af1# => X"b9050046",
		16#4af2# => X"9d080038",
		16#4af3# => X"b8680003",
		16#4af4# => X"19a00001",
		16#4af5# => X"a9adb20c",
		16#4af6# => X"e0636800",
		16#4af7# => X"84c30008",
		16#4af8# => X"e4061800",
		16#4af9# => X"10000066",
		16#4afa# => X"b9080082",
		16#4afb# => X"84e60004",
		16#4afc# => X"9d00fffc",
		16#4afd# => X"e0e74003",
		16#4afe# => X"e4853800",
		16#4aff# => X"10000009",
		16#4b00# => X"15000000",
		16#4b01# => X"0000000c",
		16#4b02# => X"8466000c",
		16#4b03# => X"84e60004",
		16#4b04# => X"e0e75803",
		16#4b05# => X"e4853800",
		16#4b06# => X"0c000006",
		16#4b07# => X"15000000",
		16#4b08# => X"84c60008",
		16#4b09# => X"e4033000",
		16#4b0a# => X"0ffffff9",
		16#4b0b# => X"9d60fffc",
		16#4b0c# => X"8466000c",
		16#4b0d# => X"d404180c",
		16#4b0e# => X"d4043008",
		16#4b0f# => X"d4032008",
		16#4b10# => X"d406200c",
		16#4b11# => X"9c21000c",
		16#4b12# => X"a8620000",
		16#4b13# => X"8521fffc",
		16#4b14# => X"8441fff4",
		16#4b15# => X"03ffe8c7",
		16#4b16# => X"85c1fff8",
		16#4b17# => X"9c21000c",
		16#4b18# => X"8521fffc",
		16#4b19# => X"8441fff4",
		16#4b1a# => X"44004800",
		16#4b1b# => X"85c1fff8",
		16#4b1c# => X"19000001",
		16#4b1d# => X"84660008",
		16#4b1e# => X"a908b214",
		16#4b1f# => X"e4234000",
		16#4b20# => X"13ffffc1",
		16#4b21# => X"15000000",
		16#4b22# => X"a8e50001",
		16#4b23# => X"e0c42800",
		16#4b24# => X"d403200c",
		16#4b25# => X"d4032008",
		16#4b26# => X"d404180c",
		16#4b27# => X"d4041808",
		16#4b28# => X"d4043804",
		16#4b29# => X"03ffffe8",
		16#4b2a# => X"d4062800",
		16#4b2b# => X"b8a50043",
		16#4b2c# => X"19600001",
		16#4b2d# => X"b8650082",
		16#4b2e# => X"b8a50003",
		16#4b2f# => X"a96bb20c",
		16#4b30# => X"e0c61808",
		16#4b31# => X"e0a55800",
		16#4b32# => X"85070004",
		16#4b33# => X"84650008",
		16#4b34# => X"e0c83004",
		16#4b35# => X"d4041808",
		16#4b36# => X"d404280c",
		16#4b37# => X"d403200c",
		16#4b38# => X"d4073004",
		16#4b39# => X"d4052008",
		16#4b3a# => X"9c21000c",
		16#4b3b# => X"a8620000",
		16#4b3c# => X"8521fffc",
		16#4b3d# => X"8441fff4",
		16#4b3e# => X"03ffe89e",
		16#4b3f# => X"85c1fff8",
		16#4b40# => X"a5080001",
		16#4b41# => X"bc280000",
		16#4b42# => X"10000009",
		16#4b43# => X"e0a32800",
		16#4b44# => X"84640000",
		16#4b45# => X"e0841802",
		16#4b46# => X"e0a51800",
		16#4b47# => X"84c40008",
		16#4b48# => X"8464000c",
		16#4b49# => X"d406180c",
		16#4b4a# => X"d4033008",
		16#4b4b# => X"a8650001",
		16#4b4c# => X"d4072008",
		16#4b4d# => X"d4041804",
		16#4b4e# => X"18600001",
		16#4b4f# => X"a863b614",
		16#4b50# => X"84630000",
		16#4b51# => X"e4851800",
		16#4b52# => X"13ffffbf",
		16#4b53# => X"18800001",
		16#4b54# => X"a8620000",
		16#4b55# => X"a884c4bc",
		16#4b56# => X"07ffff09",
		16#4b57# => X"84840000",
		16#4b58# => X"03ffffba",
		16#4b59# => X"9c21000c",
		16#4b5a# => X"1000000c",
		16#4b5b# => X"bc430054",
		16#4b5c# => X"9d03005b",
		16#4b5d# => X"03ffff97",
		16#4b5e# => X"b8680003",
		16#4b5f# => X"9c600001",
		16#4b60# => X"85670004",
		16#4b61# => X"e0a34008",
		16#4b62# => X"a8660000",
		16#4b63# => X"e0ab2804",
		16#4b64# => X"03ffffa9",
		16#4b65# => X"d4072804",
		16#4b66# => X"10000006",
		16#4b67# => X"bc430154",
		16#4b68# => X"b905004c",
		16#4b69# => X"9d08006e",
		16#4b6a# => X"03ffff8a",
		16#4b6b# => X"b8680003",
		16#4b6c# => X"10000006",
		16#4b6d# => X"bc430554",
		16#4b6e# => X"b905004f",
		16#4b6f# => X"9d080077",
		16#4b70# => X"03ffff84",
		16#4b71# => X"b8680003",
		16#4b72# => X"10000006",
		16#4b73# => X"15000000",
		16#4b74# => X"b9050052",
		16#4b75# => X"9d08007c",
		16#4b76# => X"03ffff7e",
		16#4b77# => X"b8680003",
		16#4b78# => X"9c6003f0",
		16#4b79# => X"03ffff7b",
		16#4b7a# => X"9d00007e",
		16#4b7b# => X"d7e117d4",
		16#4b7c# => X"d7e197e0",
		16#4b7d# => X"d7e1e7f4",
		16#4b7e# => X"d7e14ffc",
		16#4b7f# => X"d7e177d8",
		16#4b80# => X"d7e187dc",
		16#4b81# => X"d7e1a7e4",
		16#4b82# => X"d7e1b7e8",
		16#4b83# => X"d7e1c7ec",
		16#4b84# => X"d7e1d7f0",
		16#4b85# => X"d7e1f7f8",
		16#4b86# => X"85650008",
		16#4b87# => X"9c21ffd4",
		16#4b88# => X"aa450000",
		16#4b89# => X"ab830000",
		16#4b8a# => X"bc0b0000",
		16#4b8b# => X"10000027",
		16#4b8c# => X"a8440000",
		16#4b8d# => X"9864000c",
		16#4b8e# => X"a483ffff",
		16#4b8f# => X"a4a40008",
		16#4b90# => X"bc050000",
		16#4b91# => X"1000002e",
		16#4b92# => X"15000000",
		16#4b93# => X"84a20010",
		16#4b94# => X"bc250000",
		16#4b95# => X"0c00002a",
		16#4b96# => X"a4a40002",
		16#4b97# => X"bc050000",
		16#4b98# => X"10000033",
		16#4b99# => X"86120000",
		16#4b9a# => X"9ec00000",
		16#4b9b# => X"a9d60000",
		16#4b9c# => X"a8b60000",
		16#4b9d# => X"bc0e0000",
		16#4b9e# => X"10000067",
		16#4b9f# => X"a87c0000",
		16#4ba0# => X"a8ce0000",
		16#4ba1# => X"bcae0400",
		16#4ba2# => X"10000003",
		16#4ba3# => X"8482001c",
		16#4ba4# => X"9cc00400",
		16#4ba5# => X"85620024",
		16#4ba6# => X"48005800",
		16#4ba7# => X"15000000",
		16#4ba8# => X"bdab0000",
		16#4ba9# => X"100000c8",
		16#4baa# => X"e2d65800",
		16#4bab# => X"86920008",
		16#4bac# => X"e2945802",
		16#4bad# => X"e1ce5802",
		16#4bae# => X"bc340000",
		16#4baf# => X"13ffffed",
		16#4bb0# => X"d412a008",
		16#4bb1# => X"a9740000",
		16#4bb2# => X"9c21002c",
		16#4bb3# => X"8521fffc",
		16#4bb4# => X"8441ffd4",
		16#4bb5# => X"85c1ffd8",
		16#4bb6# => X"8601ffdc",
		16#4bb7# => X"8641ffe0",
		16#4bb8# => X"8681ffe4",
		16#4bb9# => X"86c1ffe8",
		16#4bba# => X"8701ffec",
		16#4bbb# => X"8741fff0",
		16#4bbc# => X"8781fff4",
		16#4bbd# => X"44004800",
		16#4bbe# => X"87c1fff8",
		16#4bbf# => X"a87c0000",
		16#4bc0# => X"07fff3c6",
		16#4bc1# => X"a8820000",
		16#4bc2# => X"bc2b0000",
		16#4bc3# => X"10000122",
		16#4bc4# => X"15000000",
		16#4bc5# => X"9862000c",
		16#4bc6# => X"a483ffff",
		16#4bc7# => X"a4a40002",
		16#4bc8# => X"bc050000",
		16#4bc9# => X"0fffffd1",
		16#4bca# => X"86120000",
		16#4bcb# => X"a6c40001",
		16#4bcc# => X"bc160000",
		16#4bcd# => X"1000003f",
		16#4bce# => X"a9d60000",
		16#4bcf# => X"aac50000",
		16#4bd0# => X"abc50000",
		16#4bd1# => X"ab450000",
		16#4bd2# => X"aa850000",
		16#4bd3# => X"bc140000",
		16#4bd4# => X"1000002c",
		16#4bd5# => X"bc3e0000",
		16#4bd6# => X"0c000102",
		16#4bd7# => X"a87a0000",
		16#4bd8# => X"e4b6a000",
		16#4bd9# => X"10000003",
		16#4bda# => X"ab160000",
		16#4bdb# => X"ab140000",
		16#4bdc# => X"84c20014",
		16#4bdd# => X"85c20008",
		16#4bde# => X"84620000",
		16#4bdf# => X"e1c67000",
		16#4be0# => X"e5587000",
		16#4be1# => X"10000003",
		16#4be2# => X"9c800001",
		16#4be3# => X"9c800000",
		16#4be4# => X"a48400ff",
		16#4be5# => X"bc040000",
		16#4be6# => X"0c0000db",
		16#4be7# => X"e5983000",
		16#4be8# => X"100000c5",
		16#4be9# => X"a89a0000",
		16#4bea# => X"85620024",
		16#4beb# => X"a87c0000",
		16#4bec# => X"8482001c",
		16#4bed# => X"48005800",
		16#4bee# => X"a8ba0000",
		16#4bef# => X"bdab0000",
		16#4bf0# => X"10000081",
		16#4bf1# => X"a9cb0000",
		16#4bf2# => X"e2d67002",
		16#4bf3# => X"bc360000",
		16#4bf4# => X"0c0000c6",
		16#4bf5# => X"a87c0000",
		16#4bf6# => X"85720008",
		16#4bf7# => X"e35a7000",
		16#4bf8# => X"e16b7002",
		16#4bf9# => X"e2947002",
		16#4bfa# => X"bc2b0000",
		16#4bfb# => X"0fffffb7",
		16#4bfc# => X"d4125808",
		16#4bfd# => X"bc140000",
		16#4bfe# => X"0fffffd8",
		16#4bff# => X"bc3e0000",
		16#4c00# => X"87500000",
		16#4c01# => X"86900004",
		16#4c02# => X"9fc00000",
		16#4c03# => X"03ffffd0",
		16#4c04# => X"9e100008",
		16#4c05# => X"86d00000",
		16#4c06# => X"85d00004",
		16#4c07# => X"03ffff95",
		16#4c08# => X"9e100008",
		16#4c09# => X"86d00000",
		16#4c0a# => X"85d00004",
		16#4c0b# => X"9e100008",
		16#4c0c# => X"bc0e0000",
		16#4c0d# => X"13fffffc",
		16#4c0e# => X"15000000",
		16#4c0f# => X"a463ffff",
		16#4c10# => X"a4830200",
		16#4c11# => X"bc040000",
		16#4c12# => X"10000023",
		16#4c13# => X"86820008",
		16#4c14# => X"e48ea000",
		16#4c15# => X"10000038",
		16#4c16# => X"ab540000",
		16#4c17# => X"a4830480",
		16#4c18# => X"bc240000",
		16#4c19# => X"1000005d",
		16#4c1a# => X"abd40000",
		16#4c1b# => X"84620000",
		16#4c1c# => X"aa8e0000",
		16#4c1d# => X"a8960000",
		16#4c1e# => X"a8ba0000",
		16#4c1f# => X"0400027b",
		16#4c20# => X"ab0e0000",
		16#4c21# => X"84820008",
		16#4c22# => X"84620000",
		16#4c23# => X"e3c4f002",
		16#4c24# => X"e343d000",
		16#4c25# => X"d402f008",
		16#4c26# => X"d402d000",
		16#4c27# => X"84720008",
		16#4c28# => X"e2d6c000",
		16#4c29# => X"e283a002",
		16#4c2a# => X"e1cec002",
		16#4c2b# => X"bc340000",
		16#4c2c# => X"0fffff85",
		16#4c2d# => X"d412a008",
		16#4c2e# => X"bc0e0000",
		16#4c2f# => X"0fffffe0",
		16#4c30# => X"9862000c",
		16#4c31# => X"86d00000",
		16#4c32# => X"85d00004",
		16#4c33# => X"03ffffd9",
		16#4c34# => X"9e100008",
		16#4c35# => X"84620000",
		16#4c36# => X"ab140000",
		16#4c37# => X"e4947000",
		16#4c38# => X"10000003",
		16#4c39# => X"9ca00001",
		16#4c3a# => X"a8a40000",
		16#4c3b# => X"a4a500ff",
		16#4c3c# => X"bc050000",
		16#4c3d# => X"0c000020",
		16#4c3e# => X"15000000",
		16#4c3f# => X"84c20014",
		16#4c40# => X"e48e3000",
		16#4c41# => X"10000011",
		16#4c42# => X"a8960000",
		16#4c43# => X"85620024",
		16#4c44# => X"a87c0000",
		16#4c45# => X"8482001c",
		16#4c46# => X"48005800",
		16#4c47# => X"a8b60000",
		16#4c48# => X"bdab0000",
		16#4c49# => X"10000028",
		16#4c4a# => X"aa8b0000",
		16#4c4b# => X"03ffffdc",
		16#4c4c# => X"ab0b0000",
		16#4c4d# => X"abce0000",
		16#4c4e# => X"84620000",
		16#4c4f# => X"ab4e0000",
		16#4c50# => X"03ffffcd",
		16#4c51# => X"aa8e0000",
		16#4c52# => X"a8ae0000",
		16#4c53# => X"04000247",
		16#4c54# => X"aa8e0000",
		16#4c55# => X"84820008",
		16#4c56# => X"84620000",
		16#4c57# => X"e0847002",
		16#4c58# => X"e0637000",
		16#4c59# => X"d4022008",
		16#4c5a# => X"d4021800",
		16#4c5b# => X"03ffffcc",
		16#4c5c# => X"ab0e0000",
		16#4c5d# => X"84a20010",
		16#4c5e# => X"e4432800",
		16#4c5f# => X"10000003",
		16#4c60# => X"9c800001",
		16#4c61# => X"9c800000",
		16#4c62# => X"a48400ff",
		16#4c63# => X"bc040000",
		16#4c64# => X"13ffffdb",
		16#4c65# => X"a8960000",
		16#4c66# => X"04000234",
		16#4c67# => X"a8b40000",
		16#4c68# => X"84a20000",
		16#4c69# => X"a87c0000",
		16#4c6a# => X"e0a5a000",
		16#4c6b# => X"a8820000",
		16#4c6c# => X"07fffc14",
		16#4c6d# => X"d4022800",
		16#4c6e# => X"bc2b0000",
		16#4c6f# => X"0fffffb8",
		16#4c70# => X"15000000",
		16#4c71# => X"9462000c",
		16#4c72# => X"a8630040",
		16#4c73# => X"9d60ffff",
		16#4c74# => X"03ffff3e",
		16#4c75# => X"dc02180c",
		16#4c76# => X"84a20014",
		16#4c77# => X"84820010",
		16#4c78# => X"e0c52800",
		16#4c79# => X"87420000",
		16#4c7a# => X"e0a62800",
		16#4c7b# => X"e35a2002",
		16#4c7c# => X"ba85005f",
		16#4c7d# => X"9cda0001",
		16#4c7e# => X"e0b42800",
		16#4c7f# => X"e0c67000",
		16#4c80# => X"ba850081",
		16#4c81# => X"e4743000",
		16#4c82# => X"10000004",
		16#4c83# => X"a8b40000",
		16#4c84# => X"aa860000",
		16#4c85# => X"a8a60000",
		16#4c86# => X"a4630400",
		16#4c87# => X"bc030000",
		16#4c88# => X"1000001a",
		16#4c89# => X"a87c0000",
		16#4c8a# => X"07ffe500",
		16#4c8b# => X"a8850000",
		16#4c8c# => X"bc2b0000",
		16#4c8d# => X"0c00001d",
		16#4c8e# => X"ab0b0000",
		16#4c8f# => X"a86b0000",
		16#4c90# => X"84820010",
		16#4c91# => X"040001c5",
		16#4c92# => X"a8ba0000",
		16#4c93# => X"9462000c",
		16#4c94# => X"9c80fb7f",
		16#4c95# => X"e0632003",
		16#4c96# => X"a8630080",
		16#4c97# => X"dc02180c",
		16#4c98# => X"e078d000",
		16#4c99# => X"e354d002",
		16#4c9a# => X"d402a014",
		16#4c9b# => X"d402d008",
		16#4c9c# => X"d402c010",
		16#4c9d# => X"d4021800",
		16#4c9e# => X"abce0000",
		16#4c9f# => X"ab4e0000",
		16#4ca0# => X"03ffff7d",
		16#4ca1# => X"aa8e0000",
		16#4ca2# => X"04000736",
		16#4ca3# => X"a87c0000",
		16#4ca4# => X"bc2b0000",
		16#4ca5# => X"13fffff3",
		16#4ca6# => X"ab0b0000",
		16#4ca7# => X"a87c0000",
		16#4ca8# => X"07fffe07",
		16#4ca9# => X"84820010",
		16#4caa# => X"9c60000c",
		16#4cab# => X"03ffffc6",
		16#4cac# => X"d41c1800",
		16#4cad# => X"a8b80000",
		16#4cae# => X"040001ec",
		16#4caf# => X"a9d80000",
		16#4cb0# => X"84620008",
		16#4cb1# => X"84820000",
		16#4cb2# => X"e063c002",
		16#4cb3# => X"e304c000",
		16#4cb4# => X"e2d67002",
		16#4cb5# => X"d4021808",
		16#4cb6# => X"bc360000",
		16#4cb7# => X"13ffff3f",
		16#4cb8# => X"d402c000",
		16#4cb9# => X"a87c0000",
		16#4cba# => X"07fffbc6",
		16#4cbb# => X"a8820000",
		16#4cbc# => X"bc2b0000",
		16#4cbd# => X"13ffffb4",
		16#4cbe# => X"15000000",
		16#4cbf# => X"03ffff37",
		16#4cc0# => X"abd60000",
		16#4cc1# => X"84a20010",
		16#4cc2# => X"e4432800",
		16#4cc3# => X"10000003",
		16#4cc4# => X"9c800001",
		16#4cc5# => X"9c800000",
		16#4cc6# => X"a48400ff",
		16#4cc7# => X"bc040000",
		16#4cc8# => X"13ffff20",
		16#4cc9# => X"e5983000",
		16#4cca# => X"a89a0000",
		16#4ccb# => X"040001cf",
		16#4ccc# => X"a8ae0000",
		16#4ccd# => X"84a20000",
		16#4cce# => X"a87c0000",
		16#4ccf# => X"e0a57000",
		16#4cd0# => X"a8820000",
		16#4cd1# => X"07fffbaf",
		16#4cd2# => X"d4022800",
		16#4cd3# => X"bc2b0000",
		16#4cd4# => X"0fffff1f",
		16#4cd5# => X"e2d67002",
		16#4cd6# => X"03ffff9c",
		16#4cd7# => X"9462000c",
		16#4cd8# => X"9c80000a",
		16#4cd9# => X"04000132",
		16#4cda# => X"a8b40000",
		16#4cdb# => X"bc0b0000",
		16#4cdc# => X"10000006",
		16#4cdd# => X"15000000",
		16#4cde# => X"9ecb0001",
		16#4cdf# => X"9fc00001",
		16#4ce0# => X"03fffef8",
		16#4ce1# => X"e2d6d002",
		16#4ce2# => X"9ed40001",
		16#4ce3# => X"03fffef5",
		16#4ce4# => X"9fc00001",
		16#4ce5# => X"9462000c",
		16#4ce6# => X"a8630040",
		16#4ce7# => X"9d60ffff",
		16#4ce8# => X"dc02180c",
		16#4ce9# => X"9c400009",
		16#4cea# => X"03fffec8",
		16#4ceb# => X"d41c1000",
		16#4cec# => X"d7e187f0",
		16#4ced# => X"d7e197f4",
		16#4cee# => X"d7e1a7f8",
		16#4cef# => X"d7e14ffc",
		16#4cf0# => X"d7e117e8",
		16#4cf1# => X"d7e177ec",
		16#4cf2# => X"9c21ffe8",
		16#4cf3# => X"9e0302e0",
		16#4cf4# => X"07fffd4f",
		16#4cf5# => X"aa840000",
		16#4cf6# => X"bc100000",
		16#4cf7# => X"1000001c",
		16#4cf8# => X"aa500000",
		16#4cf9# => X"9e400000",
		16#4cfa# => X"85d00004",
		16#4cfb# => X"9dceffff",
		16#4cfc# => X"bd8e0000",
		16#4cfd# => X"10000012",
		16#4cfe# => X"84500008",
		16#4cff# => X"9c42000c",
		16#4d00# => X"98620000",
		16#4d01# => X"9dceffff",
		16#4d02# => X"bc030000",
		16#4d03# => X"10000009",
		16#4d04# => X"9c62fff4",
		16#4d05# => X"98a20002",
		16#4d06# => X"bc05ffff",
		16#4d07# => X"10000006",
		16#4d08# => X"bd6e0000",
		16#4d09# => X"4800a000",
		16#4d0a# => X"15000000",
		16#4d0b# => X"e2525804",
		16#4d0c# => X"bd6e0000",
		16#4d0d# => X"13fffff3",
		16#4d0e# => X"9c420068",
		16#4d0f# => X"86100000",
		16#4d10# => X"bc300000",
		16#4d11# => X"13ffffe9",
		16#4d12# => X"15000000",
		16#4d13# => X"07fffd32",
		16#4d14# => X"15000000",
		16#4d15# => X"9c210018",
		16#4d16# => X"a9720000",
		16#4d17# => X"8521fffc",
		16#4d18# => X"8441ffe8",
		16#4d19# => X"85c1ffec",
		16#4d1a# => X"8601fff0",
		16#4d1b# => X"8641fff4",
		16#4d1c# => X"44004800",
		16#4d1d# => X"8681fff8",
		16#4d1e# => X"d7e187ec",
		16#4d1f# => X"d7e197f0",
		16#4d20# => X"d7e1a7f4",
		16#4d21# => X"d7e1b7f8",
		16#4d22# => X"d7e14ffc",
		16#4d23# => X"d7e117e4",
		16#4d24# => X"d7e177e8",
		16#4d25# => X"9c21ffe4",
		16#4d26# => X"9e0302e0",
		16#4d27# => X"aa830000",
		16#4d28# => X"07fffd1b",
		16#4d29# => X"aac40000",
		16#4d2a# => X"bc100000",
		16#4d2b# => X"1000001c",
		16#4d2c# => X"aa500000",
		16#4d2d# => X"9e400000",
		16#4d2e# => X"85d00004",
		16#4d2f# => X"9dceffff",
		16#4d30# => X"bd8e0000",
		16#4d31# => X"10000012",
		16#4d32# => X"84500008",
		16#4d33# => X"9c42000c",
		16#4d34# => X"98a20000",
		16#4d35# => X"9dceffff",
		16#4d36# => X"bc050000",
		16#4d37# => X"10000009",
		16#4d38# => X"9c82fff4",
		16#4d39# => X"98a20002",
		16#4d3a# => X"bc05ffff",
		16#4d3b# => X"10000005",
		16#4d3c# => X"a8740000",
		16#4d3d# => X"4800b000",
		16#4d3e# => X"15000000",
		16#4d3f# => X"e2525804",
		16#4d40# => X"bd6e0000",
		16#4d41# => X"13fffff3",
		16#4d42# => X"9c420068",
		16#4d43# => X"86100000",
		16#4d44# => X"bc300000",
		16#4d45# => X"13ffffe9",
		16#4d46# => X"15000000",
		16#4d47# => X"07fffcfe",
		16#4d48# => X"15000000",
		16#4d49# => X"9c21001c",
		16#4d4a# => X"a9720000",
		16#4d4b# => X"8521fffc",
		16#4d4c# => X"8441ffe4",
		16#4d4d# => X"85c1ffe8",
		16#4d4e# => X"8601ffec",
		16#4d4f# => X"8641fff0",
		16#4d50# => X"8681fff4",
		16#4d51# => X"44004800",
		16#4d52# => X"86c1fff8",
		16#4d53# => X"d7e117f4",
		16#4d54# => X"d7e177f8",
		16#4d55# => X"d7e14ffc",
		16#4d56# => X"19c00001",
		16#4d57# => X"9c21fff4",
		16#4d58# => X"a8450000",
		16#4d59# => X"bc050000",
		16#4d5a# => X"10000009",
		16#4d5b# => X"a9ce8894",
		16#4d5c# => X"18800001",
		16#4d5d# => X"a8650000",
		16#4d5e# => X"04000972",
		16#4d5f# => X"a8848abc",
		16#4d60# => X"bc0b0000",
		16#4d61# => X"0c000008",
		16#4d62# => X"a8620000",
		16#4d63# => X"9c21000c",
		16#4d64# => X"a96e0000",
		16#4d65# => X"8521fffc",
		16#4d66# => X"8441fff4",
		16#4d67# => X"44004800",
		16#4d68# => X"85c1fff8",
		16#4d69# => X"04000967",
		16#4d6a# => X"a88e0000",
		16#4d6b# => X"bc0b0000",
		16#4d6c# => X"13fffff7",
		16#4d6d# => X"a8620000",
		16#4d6e# => X"18800001",
		16#4d6f# => X"a884853b",
		16#4d70# => X"04000960",
		16#4d71# => X"9dc00000",
		16#4d72# => X"e42b7000",
		16#4d73# => X"13fffff0",
		16#4d74# => X"15000000",
		16#4d75# => X"19c00001",
		16#4d76# => X"03ffffed",
		16#4d77# => X"a9ce8894",
		16#4d78# => X"19600001",
		16#4d79# => X"44004800",
		16#4d7a# => X"a96bb7b8",
		16#4d7b# => X"19600001",
		16#4d7c# => X"44004800",
		16#4d7d# => X"a96bb798",
		16#4d7e# => X"44004800",
		16#4d7f# => X"9d600000",
		16#4d80# => X"19600001",
		16#4d81# => X"44004800",
		16#4d82# => X"a96b8ac4",
		16#4d83# => X"a8a40000",
		16#4d84# => X"a8830000",
		16#4d85# => X"18600001",
		16#4d86# => X"d7e14ffc",
		16#4d87# => X"a863ade4",
		16#4d88# => X"9c21fffc",
		16#4d89# => X"84630000",
		16#4d8a# => X"9c210004",
		16#4d8b# => X"8521fffc",
		16#4d8c# => X"03ffffc7",
		16#4d8d# => X"15000000",
		16#4d8e# => X"19600001",
		16#4d8f# => X"44004800",
		16#4d90# => X"a96b8ac4",
		16#4d91# => X"98a4000c",
		16#4d92# => X"a4c5ffff",
		16#4d93# => X"d7e117ec",
		16#4d94# => X"d7e177f0",
		16#4d95# => X"d7e14ffc",
		16#4d96# => X"d7e187f4",
		16#4d97# => X"d7e197f8",
		16#4d98# => X"a8440000",
		16#4d99# => X"a4860002",
		16#4d9a# => X"9c21ffb0",
		16#4d9b# => X"bc040000",
		16#4d9c# => X"0c000039",
		16#4d9d# => X"a9c30000",
		16#4d9e# => X"9882000e",
		16#4d9f# => X"bd840000",
		16#4da0# => X"10000018",
		16#4da1# => X"a4c60080",
		16#4da2# => X"04000f0e",
		16#4da3# => X"a8a10000",
		16#4da4# => X"bd6b0000",
		16#4da5# => X"0c000010",
		16#4da6# => X"84810004",
		16#4da7# => X"a8a08000",
		16#4da8# => X"a484f000",
		16#4da9# => X"ac642000",
		16#4daa# => X"e4242800",
		16#4dab# => X"e2401802",
		16#4dac# => X"e2521804",
		16#4dad# => X"ae52ffff",
		16#4dae# => X"0c000045",
		16#4daf# => X"ba52005f",
		16#4db0# => X"9462000c",
		16#4db1# => X"a8630800",
		16#4db2# => X"9e000400",
		16#4db3# => X"0000000b",
		16#4db4# => X"dc02180c",
		16#4db5# => X"98a2000c",
		16#4db6# => X"a4c5ffff",
		16#4db7# => X"a4c60080",
		16#4db8# => X"bc260000",
		16#4db9# => X"0c000038",
		16#4dba# => X"9e000040",
		16#4dbb# => X"a8a50800",
		16#4dbc# => X"9e400000",
		16#4dbd# => X"dc02280c",
		16#4dbe# => X"a86e0000",
		16#4dbf# => X"07ffe3cb",
		16#4dc0# => X"a8900000",
		16#4dc1# => X"bc2b0000",
		16#4dc2# => X"0c00003d",
		16#4dc3# => X"18800001",
		16#4dc4# => X"9462000c",
		16#4dc5# => X"a8630080",
		16#4dc6# => X"a8842590",
		16#4dc7# => X"bc120000",
		16#4dc8# => X"d40e203c",
		16#4dc9# => X"dc02180c",
		16#4dca# => X"d4025800",
		16#4dcb# => X"d4025810",
		16#4dcc# => X"0c000015",
		16#4dcd# => X"d4028014",
		16#4dce# => X"9c210050",
		16#4dcf# => X"8521fffc",
		16#4dd0# => X"8441ffec",
		16#4dd1# => X"85c1fff0",
		16#4dd2# => X"8601fff4",
		16#4dd3# => X"44004800",
		16#4dd4# => X"8641fff8",
		16#4dd5# => X"9c620043",
		16#4dd6# => X"d4021800",
		16#4dd7# => X"d4021810",
		16#4dd8# => X"9c600001",
		16#4dd9# => X"d4021814",
		16#4dda# => X"9c210050",
		16#4ddb# => X"8521fffc",
		16#4ddc# => X"8441ffec",
		16#4ddd# => X"85c1fff0",
		16#4dde# => X"8601fff4",
		16#4ddf# => X"44004800",
		16#4de0# => X"8641fff8",
		16#4de1# => X"9882000e",
		16#4de2# => X"04000eec",
		16#4de3# => X"a86e0000",
		16#4de4# => X"bc0b0000",
		16#4de5# => X"13ffffe9",
		16#4de6# => X"15000000",
		16#4de7# => X"9462000c",
		16#4de8# => X"a8630001",
		16#4de9# => X"dc02180c",
		16#4dea# => X"9c210050",
		16#4deb# => X"8521fffc",
		16#4dec# => X"8441ffec",
		16#4ded# => X"85c1fff0",
		16#4dee# => X"8601fff4",
		16#4def# => X"44004800",
		16#4df0# => X"8641fff8",
		16#4df1# => X"03ffffca",
		16#4df2# => X"9e000400",
		16#4df3# => X"18800001",
		16#4df4# => X"84620028",
		16#4df5# => X"a8845ac4",
		16#4df6# => X"e4232000",
		16#4df7# => X"13ffffb9",
		16#4df8# => X"15000000",
		16#4df9# => X"9462000c",
		16#4dfa# => X"9e000400",
		16#4dfb# => X"e0638004",
		16#4dfc# => X"d402804c",
		16#4dfd# => X"03ffffc1",
		16#4dfe# => X"dc02180c",
		16#4dff# => X"9862000c",
		16#4e00# => X"a4830200",
		16#4e01# => X"bc240000",
		16#4e02# => X"13ffffcc",
		16#4e03# => X"a8630002",
		16#4e04# => X"9c820043",
		16#4e05# => X"dc02180c",
		16#4e06# => X"9c600001",
		16#4e07# => X"d4022000",
		16#4e08# => X"d4022010",
		16#4e09# => X"03ffffc5",
		16#4e0a# => X"d4021814",
		16#4e0b# => X"d7e117fc",
		16#4e0c# => X"a4c30003",
		16#4e0d# => X"9c21fffc",
		16#4e0e# => X"bc060000",
		16#4e0f# => X"10000016",
		16#4e10# => X"a48400ff",
		16#4e11# => X"bc050000",
		16#4e12# => X"10000027",
		16#4e13# => X"a9650000",
		16#4e14# => X"8cc30000",
		16#4e15# => X"e4062000",
		16#4e16# => X"10000023",
		16#4e17# => X"a9630000",
		16#4e18# => X"00000008",
		16#4e19# => X"9ca5ffff",
		16#4e1a# => X"1000001f",
		16#4e1b# => X"a9650000",
		16#4e1c# => X"8cc30000",
		16#4e1d# => X"e4062000",
		16#4e1e# => X"1000001e",
		16#4e1f# => X"9ca5ffff",
		16#4e20# => X"9c630001",
		16#4e21# => X"a4c30003",
		16#4e22# => X"bc260000",
		16#4e23# => X"13fffff7",
		16#4e24# => X"bc050000",
		16#4e25# => X"bca50003",
		16#4e26# => X"0c00001a",
		16#4e27# => X"b8c40008",
		16#4e28# => X"bc050000",
		16#4e29# => X"10000010",
		16#4e2a# => X"a9650000",
		16#4e2b# => X"8cc30000",
		16#4e2c# => X"e4062000",
		16#4e2d# => X"1000000c",
		16#4e2e# => X"a9630000",
		16#4e2f# => X"00000006",
		16#4e30# => X"9ca5ffff",
		16#4e31# => X"8cc30000",
		16#4e32# => X"e4062000",
		16#4e33# => X"10000009",
		16#4e34# => X"9ca5ffff",
		16#4e35# => X"bc250000",
		16#4e36# => X"13fffffb",
		16#4e37# => X"9c630001",
		16#4e38# => X"a9650000",
		16#4e39# => X"9c210004",
		16#4e3a# => X"44004800",
		16#4e3b# => X"8441fffc",
		16#4e3c# => X"9c210004",
		16#4e3d# => X"a9630000",
		16#4e3e# => X"44004800",
		16#4e3f# => X"8441fffc",
		16#4e40# => X"e0c62004",
		16#4e41# => X"b9060010",
		16#4e42# => X"e1083004",
		16#4e43# => X"84c30000",
		16#4e44# => X"1840fefe",
		16#4e45# => X"e0c83005",
		16#4e46# => X"a842feff",
		16#4e47# => X"e0e61000",
		16#4e48# => X"acc6ffff",
		16#4e49# => X"18408080",
		16#4e4a# => X"e0c73003",
		16#4e4b# => X"a8428080",
		16#4e4c# => X"e0c61003",
		16#4e4d# => X"bc260000",
		16#4e4e# => X"13ffffdb",
		16#4e4f# => X"bc050000",
		16#4e50# => X"9ca5fffc",
		16#4e51# => X"bc450003",
		16#4e52# => X"13fffff1",
		16#4e53# => X"9c630004",
		16#4e54# => X"03ffffd5",
		16#4e55# => X"bc050000",
		16#4e56# => X"a9030000",
		16#4e57# => X"a9840000",
		16#4e58# => X"bca5000f",
		16#4e59# => X"10000007",
		16#4e5a# => X"a8e50000",
		16#4e5b# => X"e0c41804",
		16#4e5c# => X"a4c60003",
		16#4e5d# => X"bc260000",
		16#4e5e# => X"0c00000f",
		16#4e5f# => X"a8c40000",
		16#4e60# => X"bc070000",
		16#4e61# => X"1000000a",
		16#4e62# => X"15000000",
		16#4e63# => X"9c800000",
		16#4e64# => X"e0cc2000",
		16#4e65# => X"e0a82000",
		16#4e66# => X"8cc60000",
		16#4e67# => X"9c840001",
		16#4e68# => X"e4243800",
		16#4e69# => X"13fffffb",
		16#4e6a# => X"d8053000",
		16#4e6b# => X"44004800",
		16#4e6c# => X"a9630000",
		16#4e6d# => X"a9050000",
		16#4e6e# => X"a8e30000",
		16#4e6f# => X"85660000",
		16#4e70# => X"9d08fff0",
		16#4e71# => X"d4075800",
		16#4e72# => X"bc48000f",
		16#4e73# => X"85660004",
		16#4e74# => X"d4075804",
		16#4e75# => X"85660008",
		16#4e76# => X"d4075808",
		16#4e77# => X"8566000c",
		16#4e78# => X"9cc60010",
		16#4e79# => X"d407580c",
		16#4e7a# => X"13fffff5",
		16#4e7b# => X"9ce70010",
		16#4e7c# => X"9ca5fff0",
		16#4e7d# => X"b8c50044",
		16#4e7e# => X"9d860001",
		16#4e7f# => X"b8c60004",
		16#4e80# => X"b98c0004",
		16#4e81# => X"e0a53002",
		16#4e82# => X"e1036000",
		16#4e83# => X"a8e50000",
		16#4e84# => X"bca50003",
		16#4e85# => X"13ffffdb",
		16#4e86# => X"e1846000",
		16#4e87# => X"9c800000",
		16#4e88# => X"e0cc2000",
		16#4e89# => X"e0e82000",
		16#4e8a# => X"84c60000",
		16#4e8b# => X"9c840004",
		16#4e8c# => X"d4073000",
		16#4e8d# => X"e0c52002",
		16#4e8e# => X"bc460003",
		16#4e8f# => X"13fffffa",
		16#4e90# => X"e0cc2000",
		16#4e91# => X"9ca5fffc",
		16#4e92# => X"b8e50042",
		16#4e93# => X"9c870001",
		16#4e94# => X"b8e70002",
		16#4e95# => X"b8840002",
		16#4e96# => X"e0e53802",
		16#4e97# => X"e1082000",
		16#4e98# => X"03ffffc8",
		16#4e99# => X"e18c2000",
		16#4e9a# => X"d7e117fc",
		16#4e9b# => X"a9030000",
		16#4e9c# => X"9c21fffc",
		16#4e9d# => X"a9640000",
		16#4e9e# => X"e4a32000",
		16#4e9f# => X"10000016",
		16#4ea0# => X"a8e50000",
		16#4ea1# => X"e0c42800",
		16#4ea2# => X"e4633000",
		16#4ea3# => X"10000013",
		16#4ea4# => X"bca5000f",
		16#4ea5# => X"bc050000",
		16#4ea6# => X"1000000b",
		16#4ea7# => X"15000000",
		16#4ea8# => X"e0832800",
		16#4ea9# => X"9ca5ffff",
		16#4eaa# => X"9cc6ffff",
		16#4eab# => X"9c84ffff",
		16#4eac# => X"8c460000",
		16#4ead# => X"9ca5ffff",
		16#4eae# => X"bc25ffff",
		16#4eaf# => X"13fffffb",
		16#4eb0# => X"d8041000",
		16#4eb1# => X"9c210004",
		16#4eb2# => X"a9630000",
		16#4eb3# => X"44004800",
		16#4eb4# => X"8441fffc",
		16#4eb5# => X"bca5000f",
		16#4eb6# => X"0c000011",
		16#4eb7# => X"e0c41804",
		16#4eb8# => X"bc070000",
		16#4eb9# => X"13fffff8",
		16#4eba# => X"15000000",
		16#4ebb# => X"9c800000",
		16#4ebc# => X"e0cb2000",
		16#4ebd# => X"e0a82000",
		16#4ebe# => X"8cc60000",
		16#4ebf# => X"9c840001",
		16#4ec0# => X"e4243800",
		16#4ec1# => X"13fffffb",
		16#4ec2# => X"d8053000",
		16#4ec3# => X"9c210004",
		16#4ec4# => X"a9630000",
		16#4ec5# => X"44004800",
		16#4ec6# => X"8441fffc",
		16#4ec7# => X"a4c60003",
		16#4ec8# => X"bc260000",
		16#4ec9# => X"13fffff0",
		16#4eca# => X"bc070000",
		16#4ecb# => X"a9050000",
		16#4ecc# => X"a8c40000",
		16#4ecd# => X"a8e30000",
		16#4ece# => X"85660000",
		16#4ecf# => X"9d08fff0",
		16#4ed0# => X"d4075800",
		16#4ed1# => X"bc48000f",
		16#4ed2# => X"85660004",
		16#4ed3# => X"d4075804",
		16#4ed4# => X"85660008",
		16#4ed5# => X"d4075808",
		16#4ed6# => X"8566000c",
		16#4ed7# => X"9cc60010",
		16#4ed8# => X"d407580c",
		16#4ed9# => X"13fffff5",
		16#4eda# => X"9ce70010",
		16#4edb# => X"9ca5fff0",
		16#4edc# => X"b8c50044",
		16#4edd# => X"9d660001",
		16#4ede# => X"b8c60004",
		16#4edf# => X"b96b0004",
		16#4ee0# => X"e0a53002",
		16#4ee1# => X"e1035800",
		16#4ee2# => X"a8e50000",
		16#4ee3# => X"bca50003",
		16#4ee4# => X"13ffffd4",
		16#4ee5# => X"e1645800",
		16#4ee6# => X"9c800000",
		16#4ee7# => X"e0cb2000",
		16#4ee8# => X"e0e82000",
		16#4ee9# => X"84c60000",
		16#4eea# => X"9c840004",
		16#4eeb# => X"d4073000",
		16#4eec# => X"e0c52002",
		16#4eed# => X"bc460003",
		16#4eee# => X"13fffffa",
		16#4eef# => X"e0cb2000",
		16#4ef0# => X"9ca5fffc",
		16#4ef1# => X"b8e50042",
		16#4ef2# => X"9c870001",
		16#4ef3# => X"b8e70002",
		16#4ef4# => X"b8840002",
		16#4ef5# => X"e0e53802",
		16#4ef6# => X"e1082000",
		16#4ef7# => X"03ffffc1",
		16#4ef8# => X"e16b2000",
		16#4ef9# => X"d7e117fc",
		16#4efa# => X"a4e30003",
		16#4efb# => X"9c21fffc",
		16#4efc# => X"bc070000",
		16#4efd# => X"10000011",
		16#4efe# => X"a8c30000",
		16#4eff# => X"bc050000",
		16#4f00# => X"10000045",
		16#4f01# => X"15000000",
		16#4f02# => X"b9040018",
		16#4f03# => X"9ca5ffff",
		16#4f04# => X"00000004",
		16#4f05# => X"b9080098",
		16#4f06# => X"1000003f",
		16#4f07# => X"9ca5ffff",
		16#4f08# => X"d8064000",
		16#4f09# => X"9cc60001",
		16#4f0a# => X"a4e60003",
		16#4f0b# => X"bc270000",
		16#4f0c# => X"13fffffa",
		16#4f0d# => X"bc050000",
		16#4f0e# => X"bca50003",
		16#4f0f# => X"1000002c",
		16#4f10# => X"bc050000",
		16#4f11# => X"a50400ff",
		16#4f12# => X"a8e60000",
		16#4f13# => X"b9680008",
		16#4f14# => X"bc45000f",
		16#4f15# => X"e10b4004",
		16#4f16# => X"b9680010",
		16#4f17# => X"0c000014",
		16#4f18# => X"e10b4004",
		16#4f19# => X"a8e60000",
		16#4f1a# => X"a9850000",
		16#4f1b# => X"d4074000",
		16#4f1c# => X"d4074004",
		16#4f1d# => X"d4074008",
		16#4f1e# => X"d407400c",
		16#4f1f# => X"9d8cfff0",
		16#4f20# => X"bc4c000f",
		16#4f21# => X"13fffffa",
		16#4f22# => X"9ce70010",
		16#4f23# => X"9ca5fff0",
		16#4f24# => X"9c40fff0",
		16#4f25# => X"e0e51003",
		16#4f26# => X"a4a5000f",
		16#4f27# => X"9ce70010",
		16#4f28# => X"bc450003",
		16#4f29# => X"0c000010",
		16#4f2a# => X"e0e63800",
		16#4f2b# => X"9cc00000",
		16#4f2c# => X"e1673000",
		16#4f2d# => X"9cc60004",
		16#4f2e# => X"d40b4000",
		16#4f2f# => X"e1653002",
		16#4f30# => X"bc4b0003",
		16#4f31# => X"13fffffc",
		16#4f32# => X"e1673000",
		16#4f33# => X"9ca5fffc",
		16#4f34# => X"9c40fffc",
		16#4f35# => X"e0c51003",
		16#4f36# => X"a4a50003",
		16#4f37# => X"9cc60004",
		16#4f38# => X"e0e73000",
		16#4f39# => X"a8c70000",
		16#4f3a# => X"bc050000",
		16#4f3b# => X"1000000a",
		16#4f3c# => X"15000000",
		16#4f3d# => X"b8840018",
		16#4f3e# => X"9ce00000",
		16#4f3f# => X"b9040098",
		16#4f40# => X"e0863800",
		16#4f41# => X"9ce70001",
		16#4f42# => X"e4253800",
		16#4f43# => X"13fffffd",
		16#4f44# => X"d8044000",
		16#4f45# => X"9c210004",
		16#4f46# => X"a9630000",
		16#4f47# => X"44004800",
		16#4f48# => X"8441fffc",
		16#4f49# => X"d7e117f4",
		16#4f4a# => X"d7e177f8",
		16#4f4b# => X"d7e14ffc",
		16#4f4c# => X"a8440000",
		16#4f4d# => X"8483004c",
		16#4f4e# => X"9c21fff4",
		16#4f4f# => X"bc240000",
		16#4f50# => X"0c000012",
		16#4f51# => X"a9c30000",
		16#4f52# => X"b8620002",
		16#4f53# => X"e0841800",
		16#4f54# => X"85640000",
		16#4f55# => X"bc0b0000",
		16#4f56# => X"10000015",
		16#4f57# => X"a86e0000",
		16#4f58# => X"844b0000",
		16#4f59# => X"d4041000",
		16#4f5a# => X"9c400000",
		16#4f5b# => X"d40b1010",
		16#4f5c# => X"d40b100c",
		16#4f5d# => X"9c21000c",
		16#4f5e# => X"8521fffc",
		16#4f5f# => X"8441fff4",
		16#4f60# => X"44004800",
		16#4f61# => X"85c1fff8",
		16#4f62# => X"9c800004",
		16#4f63# => X"04000c14",
		16#4f64# => X"9ca00021",
		16#4f65# => X"a88b0000",
		16#4f66# => X"bc040000",
		16#4f67# => X"0fffffeb",
		16#4f68# => X"d40e584c",
		16#4f69# => X"03fffff5",
		16#4f6a# => X"9c21000c",
		16#4f6b# => X"9c800001",
		16#4f6c# => X"e1c41008",
		16#4f6d# => X"9cae0005",
		16#4f6e# => X"04000c09",
		16#4f6f# => X"b8a50002",
		16#4f70# => X"bc0b0000",
		16#4f71# => X"13ffffec",
		16#4f72# => X"15000000",
		16#4f73# => X"d40b1004",
		16#4f74# => X"03ffffe6",
		16#4f75# => X"d40b7008",
		16#4f76# => X"bc040000",
		16#4f77# => X"10000009",
		16#4f78# => X"15000000",
		16#4f79# => X"84c40004",
		16#4f7a# => X"84a3004c",
		16#4f7b# => X"b8660002",
		16#4f7c# => X"e0651800",
		16#4f7d# => X"84a30000",
		16#4f7e# => X"d4042800",
		16#4f7f# => X"d4032000",
		16#4f80# => X"44004800",
		16#4f81# => X"15000000",
		16#4f82# => X"d7e117e8",
		16#4f83# => X"d7e177ec",
		16#4f84# => X"d7e187f0",
		16#4f85# => X"d7e197f4",
		16#4f86# => X"d7e14ffc",
		16#4f87# => X"d7e1a7f8",
		16#4f88# => X"a9c40000",
		16#4f89# => X"9c21ffe8",
		16#4f8a# => X"aa430000",
		16#4f8b# => X"a8460000",
		16#4f8c# => X"86040010",
		16#4f8d# => X"9ce40014",
		16#4f8e# => X"9d000000",
		16#4f8f# => X"84870000",
		16#4f90# => X"9d080001",
		16#4f91# => X"a4c4ffff",
		16#4f92# => X"b8840050",
		16#4f93# => X"e0c53306",
		16#4f94# => X"e0852306",
		16#4f95# => X"e0c23000",
		16#4f96# => X"e5504000",
		16#4f97# => X"b8460050",
		16#4f98# => X"a4c6ffff",
		16#4f99# => X"e0422000",
		16#4f9a# => X"b8820010",
		16#4f9b# => X"b8420050",
		16#4f9c# => X"e0c43000",
		16#4f9d# => X"d4073000",
		16#4f9e# => X"13fffff1",
		16#4f9f# => X"9ce70004",
		16#4fa0# => X"bc020000",
		16#4fa1# => X"1000000c",
		16#4fa2# => X"15000000",
		16#4fa3# => X"846e0008",
		16#4fa4# => X"e5901800",
		16#4fa5# => X"0c000011",
		16#4fa6# => X"a8720000",
		16#4fa7# => X"9c700005",
		16#4fa8# => X"9e100001",
		16#4fa9# => X"b8630002",
		16#4faa# => X"d40e8010",
		16#4fab# => X"e06e1800",
		16#4fac# => X"d4031000",
		16#4fad# => X"9c210018",
		16#4fae# => X"a96e0000",
		16#4faf# => X"8521fffc",
		16#4fb0# => X"8441ffe8",
		16#4fb1# => X"85c1ffec",
		16#4fb2# => X"8601fff0",
		16#4fb3# => X"8641fff4",
		16#4fb4# => X"44004800",
		16#4fb5# => X"8681fff8",
		16#4fb6# => X"848e0004",
		16#4fb7# => X"07ffff92",
		16#4fb8# => X"9c840001",
		16#4fb9# => X"84ae0010",
		16#4fba# => X"9c8e000c",
		16#4fbb# => X"9ca50002",
		16#4fbc# => X"9c6b000c",
		16#4fbd# => X"b8a50002",
		16#4fbe# => X"07fffe98",
		16#4fbf# => X"aa8b0000",
		16#4fc0# => X"846e0004",
		16#4fc1# => X"8492004c",
		16#4fc2# => X"b8630002",
		16#4fc3# => X"e0641800",
		16#4fc4# => X"84830000",
		16#4fc5# => X"d40e2000",
		16#4fc6# => X"d4037000",
		16#4fc7# => X"03ffffe0",
		16#4fc8# => X"a9d40000",
		16#4fc9# => X"d7e177e8",
		16#4fca# => X"d7e187ec",
		16#4fcb# => X"d7e197f0",
		16#4fcc# => X"d7e1a7f4",
		16#4fcd# => X"d7e1b7f8",
		16#4fce# => X"d7e14ffc",
		16#4fcf# => X"d7e117e4",
		16#4fd0# => X"a9c30000",
		16#4fd1# => X"9c21ffe4",
		16#4fd2# => X"aa840000",
		16#4fd3# => X"9c660008",
		16#4fd4# => X"9c800009",
		16#4fd5# => X"aa060000",
		16#4fd6# => X"aa450000",
		16#4fd7# => X"07ffd634",
		16#4fd8# => X"aac70000",
		16#4fd9# => X"bdab0001",
		16#4fda# => X"10000007",
		16#4fdb# => X"9c800000",
		16#4fdc# => X"9c400001",
		16#4fdd# => X"e0421000",
		16#4fde# => X"e54b1000",
		16#4fdf# => X"13fffffe",
		16#4fe0# => X"9c840001",
		16#4fe1# => X"a86e0000",
		16#4fe2# => X"07ffff67",
		16#4fe3# => X"9c400001",
		16#4fe4# => X"d40bb014",
		16#4fe5# => X"bdb20009",
		16#4fe6# => X"10000029",
		16#4fe7# => X"d40b1010",
		16#4fe8# => X"9ed40009",
		16#4fe9# => X"9c400009",
		16#4fea# => X"e0941000",
		16#4feb# => X"a86e0000",
		16#4fec# => X"90c40000",
		16#4fed# => X"9ca0000a",
		16#4fee# => X"a88b0000",
		16#4fef# => X"9cc6ffd0",
		16#4ff0# => X"07ffff92",
		16#4ff1# => X"9c420001",
		16#4ff2# => X"e5521000",
		16#4ff3# => X"13fffff8",
		16#4ff4# => X"e0941000",
		16#4ff5# => X"e2969000",
		16#4ff6# => X"9e94fff8",
		16#4ff7# => X"e5b09000",
		16#4ff8# => X"1000000e",
		16#4ff9# => X"9c400000",
		16#4ffa# => X"e0941000",
		16#4ffb# => X"a86e0000",
		16#4ffc# => X"90e40000",
		16#4ffd# => X"9ca0000a",
		16#4ffe# => X"a88b0000",
		16#4fff# => X"9cc7ffd0",
		16#5000# => X"07ffff82",
		16#5001# => X"9c420001",
		16#5002# => X"e0629000",
		16#5003# => X"e5501800",
		16#5004# => X"13fffff7",
		16#5005# => X"e0941000",
		16#5006# => X"9c21001c",
		16#5007# => X"8521fffc",
		16#5008# => X"8441ffe4",
		16#5009# => X"85c1ffe8",
		16#500a# => X"8601ffec",
		16#500b# => X"8641fff0",
		16#500c# => X"8681fff4",
		16#500d# => X"44004800",
		16#500e# => X"86c1fff8",
		16#500f# => X"9e94000a",
		16#5010# => X"03ffffe7",
		16#5011# => X"9e400009",
		16#5012# => X"d7e117fc",
		16#5013# => X"1840ffff",
		16#5014# => X"9d600000",
		16#5015# => X"e0831003",
		16#5016# => X"e4245800",
		16#5017# => X"10000004",
		16#5018# => X"9c21fffc",
		16#5019# => X"b8630010",
		16#501a# => X"9d600010",
		16#501b# => X"1840ff00",
		16#501c# => X"e0831003",
		16#501d# => X"bc240000",
		16#501e# => X"10000004",
		16#501f# => X"1840f000",
		16#5020# => X"b8630008",
		16#5021# => X"9d6b0008",
		16#5022# => X"e0831003",
		16#5023# => X"bc240000",
		16#5024# => X"10000004",
		16#5025# => X"1840c000",
		16#5026# => X"b8630004",
		16#5027# => X"9d6b0004",
		16#5028# => X"e0831003",
		16#5029# => X"bc240000",
		16#502a# => X"10000005",
		16#502b# => X"bd830000",
		16#502c# => X"b8630002",
		16#502d# => X"9d6b0002",
		16#502e# => X"bd830000",
		16#502f# => X"10000007",
		16#5030# => X"15000000",
		16#5031# => X"18404000",
		16#5032# => X"e0631003",
		16#5033# => X"bc030000",
		16#5034# => X"10000005",
		16#5035# => X"9d6b0001",
		16#5036# => X"9c210004",
		16#5037# => X"44004800",
		16#5038# => X"8441fffc",
		16#5039# => X"9c210004",
		16#503a# => X"9d600020",
		16#503b# => X"44004800",
		16#503c# => X"8441fffc",
		16#503d# => X"84830000",
		16#503e# => X"a5640007",
		16#503f# => X"bc0b0000",
		16#5040# => X"1000000e",
		16#5041# => X"a4a4ffff",
		16#5042# => X"a4a40001",
		16#5043# => X"9d600000",
		16#5044# => X"e4255800",
		16#5045# => X"10000007",
		16#5046# => X"a4a40002",
		16#5047# => X"e4055800",
		16#5048# => X"0c00002a",
		16#5049# => X"9d600002",
		16#504a# => X"b8840042",
		16#504b# => X"d4032000",
		16#504c# => X"44004800",
		16#504d# => X"15000000",
		16#504e# => X"bc250000",
		16#504f# => X"10000005",
		16#5050# => X"a4a400ff",
		16#5051# => X"b8840050",
		16#5052# => X"9d600010",
		16#5053# => X"a4a400ff",
		16#5054# => X"bc250000",
		16#5055# => X"10000005",
		16#5056# => X"a4a4000f",
		16#5057# => X"b8840048",
		16#5058# => X"9d6b0008",
		16#5059# => X"a4a4000f",
		16#505a# => X"bc250000",
		16#505b# => X"10000005",
		16#505c# => X"a4a40003",
		16#505d# => X"b8840044",
		16#505e# => X"9d6b0004",
		16#505f# => X"a4a40003",
		16#5060# => X"bc250000",
		16#5061# => X"10000005",
		16#5062# => X"a4a40001",
		16#5063# => X"b8840042",
		16#5064# => X"9d6b0002",
		16#5065# => X"a4a40001",
		16#5066# => X"bc250000",
		16#5067# => X"10000007",
		16#5068# => X"15000000",
		16#5069# => X"b8840041",
		16#506a# => X"bc040000",
		16#506b# => X"10000005",
		16#506c# => X"15000000",
		16#506d# => X"9d6b0001",
		16#506e# => X"44004800",
		16#506f# => X"d4032000",
		16#5070# => X"44004800",
		16#5071# => X"9d600020",
		16#5072# => X"b8840041",
		16#5073# => X"9d600001",
		16#5074# => X"44004800",
		16#5075# => X"d4032000",
		16#5076# => X"d7e14ffc",
		16#5077# => X"d7e117f8",
		16#5078# => X"a8440000",
		16#5079# => X"9c21fff8",
		16#507a# => X"07fffecf",
		16#507b# => X"9c800001",
		16#507c# => X"9c800001",
		16#507d# => X"d40b1014",
		16#507e# => X"d40b2010",
		16#507f# => X"9c210008",
		16#5080# => X"8521fffc",
		16#5081# => X"44004800",
		16#5082# => X"8441fff8",
		16#5083# => X"d7e177ec",
		16#5084# => X"d7e187f0",
		16#5085# => X"d7e197f4",
		16#5086# => X"d7e1a7f8",
		16#5087# => X"d7e14ffc",
		16#5088# => X"d7e117e8",
		16#5089# => X"86440010",
		16#508a# => X"86850010",
		16#508b# => X"9c21ffe8",
		16#508c# => X"a9c40000",
		16#508d# => X"e572a000",
		16#508e# => X"10000008",
		16#508f# => X"aa050000",
		16#5090# => X"a8920000",
		16#5091# => X"a84e0000",
		16#5092# => X"aa540000",
		16#5093# => X"a9c50000",
		16#5094# => X"aa840000",
		16#5095# => X"aa020000",
		16#5096# => X"e0549000",
		16#5097# => X"84ae0008",
		16#5098# => X"e5a22800",
		16#5099# => X"10000003",
		16#509a# => X"848e0004",
		16#509b# => X"9c840001",
		16#509c# => X"07fffead",
		16#509d# => X"15000000",
		16#509e# => X"9ea20005",
		16#509f# => X"9e6b0014",
		16#50a0# => X"bab50002",
		16#50a1# => X"e2aba800",
		16#50a2# => X"e473a800",
		16#50a3# => X"10000009",
		16#50a4# => X"9ef40005",
		16#50a5# => X"a8d30000",
		16#50a6# => X"9c600000",
		16#50a7# => X"d4061800",
		16#50a8# => X"9cc60004",
		16#50a9# => X"e4553000",
		16#50aa# => X"13fffffd",
		16#50ab# => X"9ef40005",
		16#50ac# => X"9d920005",
		16#50ad# => X"baf70002",
		16#50ae# => X"b98c0002",
		16#50af# => X"9e300014",
		16#50b0# => X"e2f0b800",
		16#50b1# => X"9f2e0014",
		16#50b2# => X"e471b800",
		16#50b3# => X"10000045",
		16#50b4# => X"e18e6000",
		16#50b5# => X"84f10000",
		16#50b6# => X"a4a7ffff",
		16#50b7# => X"bc050000",
		16#50b8# => X"1000001e",
		16#50b9# => X"b8e70050",
		16#50ba# => X"a8730000",
		16#50bb# => X"a8990000",
		16#50bc# => X"9cc00000",
		16#50bd# => X"85a40000",
		16#50be# => X"85030000",
		16#50bf# => X"a4edffff",
		16#50c0# => X"b9ad0050",
		16#50c1# => X"e0e72b06",
		16#50c2# => X"e1ad2b06",
		16#50c3# => X"a5e8ffff",
		16#50c4# => X"b9080050",
		16#50c5# => X"e0e77800",
		16#50c6# => X"9c840004",
		16#50c7# => X"e0e73000",
		16#50c8# => X"e0cd4000",
		16#50c9# => X"b9070050",
		16#50ca# => X"a4e7ffff",
		16#50cb# => X"e44c2000",
		16#50cc# => X"e0c64000",
		16#50cd# => X"b9060010",
		16#50ce# => X"b8c60050",
		16#50cf# => X"e0e83804",
		16#50d0# => X"d4033800",
		16#50d1# => X"13ffffec",
		16#50d2# => X"9c630004",
		16#50d3# => X"d4033000",
		16#50d4# => X"84f10000",
		16#50d5# => X"b8e70050",
		16#50d6# => X"bc070000",
		16#50d7# => X"1000001d",
		16#50d8# => X"a8930000",
		16#50d9# => X"84b30000",
		16#50da# => X"a8c50000",
		16#50db# => X"a8790000",
		16#50dc# => X"9d000000",
		16#50dd# => X"85a30000",
		16#50de# => X"b8c60050",
		16#50df# => X"a5adffff",
		16#50e0# => X"a4a5ffff",
		16#50e1# => X"e1a76b06",
		16#50e2# => X"e1086800",
		16#50e3# => X"e0c83000",
		16#50e4# => X"b9a60010",
		16#50e5# => X"b9060050",
		16#50e6# => X"e0ad2804",
		16#50e7# => X"d4042800",
		16#50e8# => X"9c840004",
		16#50e9# => X"94a30000",
		16#50ea# => X"e0a72b06",
		16#50eb# => X"84c40000",
		16#50ec# => X"9c630004",
		16#50ed# => X"a5a6ffff",
		16#50ee# => X"e44c1800",
		16#50ef# => X"e0a56800",
		16#50f0# => X"e0a54000",
		16#50f1# => X"13ffffec",
		16#50f2# => X"b9050050",
		16#50f3# => X"d4042800",
		16#50f4# => X"9e310004",
		16#50f5# => X"e4b78800",
		16#50f6# => X"0fffffbf",
		16#50f7# => X"9e730004",
		16#50f8# => X"bda20000",
		16#50f9# => X"10000012",
		16#50fa# => X"15000000",
		16#50fb# => X"9c75fffc",
		16#50fc# => X"84830000",
		16#50fd# => X"bc240000",
		16#50fe# => X"0c00000a",
		16#50ff# => X"9c42ffff",
		16#5100# => X"9c420001",
		16#5101# => X"0000000b",
		16#5102# => X"d40b1010",
		16#5103# => X"84830000",
		16#5104# => X"bc040000",
		16#5105# => X"0c000006",
		16#5106# => X"15000000",
		16#5107# => X"9c42ffff",
		16#5108# => X"bda20000",
		16#5109# => X"0ffffffa",
		16#510a# => X"9c63fffc",
		16#510b# => X"d40b1010",
		16#510c# => X"9c210018",
		16#510d# => X"8521fffc",
		16#510e# => X"8441ffe8",
		16#510f# => X"85c1ffec",
		16#5110# => X"8601fff0",
		16#5111# => X"8641fff4",
		16#5112# => X"44004800",
		16#5113# => X"8681fff8",
		16#5114# => X"d7e117e8",
		16#5115# => X"d7e187f0",
		16#5116# => X"d7e1a7f8",
		16#5117# => X"d7e14ffc",
		16#5118# => X"d7e177ec",
		16#5119# => X"d7e197f4",
		16#511a# => X"a8450000",
		16#511b# => X"a4a50003",
		16#511c# => X"9c21ffe8",
		16#511d# => X"aa830000",
		16#511e# => X"bc050000",
		16#511f# => X"0c00003c",
		16#5120# => X"aa040000",
		16#5121# => X"b8420082",
		16#5122# => X"bc020000",
		16#5123# => X"10000026",
		16#5124# => X"15000000",
		16#5125# => X"85d40048",
		16#5126# => X"bc2e0000",
		16#5127# => X"1000000e",
		16#5128# => X"a4820001",
		16#5129# => X"0000003c",
		16#512a# => X"a8740000",
		16#512b# => X"b8420081",
		16#512c# => X"bc020000",
		16#512d# => X"1000001c",
		16#512e# => X"15000000",
		16#512f# => X"864e0000",
		16#5130# => X"bc320000",
		16#5131# => X"0c000021",
		16#5132# => X"a88e0000",
		16#5133# => X"a9d20000",
		16#5134# => X"a4820001",
		16#5135# => X"bc040000",
		16#5136# => X"13fffff5",
		16#5137# => X"a8900000",
		16#5138# => X"a8ae0000",
		16#5139# => X"07ffff4a",
		16#513a# => X"a8740000",
		16#513b# => X"bc100000",
		16#513c# => X"1000001d",
		16#513d# => X"15000000",
		16#513e# => X"84700004",
		16#513f# => X"8494004c",
		16#5140# => X"b8630002",
		16#5141# => X"b8420081",
		16#5142# => X"e0641800",
		16#5143# => X"bc020000",
		16#5144# => X"84830000",
		16#5145# => X"d4102000",
		16#5146# => X"d4038000",
		16#5147# => X"0fffffe8",
		16#5148# => X"aa0b0000",
		16#5149# => X"9c210018",
		16#514a# => X"a9700000",
		16#514b# => X"8521fffc",
		16#514c# => X"8441ffe8",
		16#514d# => X"85c1ffec",
		16#514e# => X"8601fff0",
		16#514f# => X"8641fff4",
		16#5150# => X"44004800",
		16#5151# => X"8681fff8",
		16#5152# => X"a8ae0000",
		16#5153# => X"07ffff30",
		16#5154# => X"a8740000",
		16#5155# => X"d40e5800",
		16#5156# => X"d40b9000",
		16#5157# => X"03ffffdd",
		16#5158# => X"a9cb0000",
		16#5159# => X"03ffffd2",
		16#515a# => X"aa0b0000",
		16#515b# => X"9ca5ffff",
		16#515c# => X"18e00001",
		16#515d# => X"b8a50002",
		16#515e# => X"a8e78c1c",
		16#515f# => X"9cc00000",
		16#5160# => X"e0a53800",
		16#5161# => X"07fffe21",
		16#5162# => X"84a50000",
		16#5163# => X"03ffffbe",
		16#5164# => X"aa0b0000",
		16#5165# => X"07ffff11",
		16#5166# => X"9c800271",
		16#5167# => X"9c600000",
		16#5168# => X"d4145848",
		16#5169# => X"a9cb0000",
		16#516a# => X"03ffffca",
		16#516b# => X"d40b1800",
		16#516c# => X"d7e177ec",
		16#516d# => X"85c40010",
		16#516e# => X"d7e187f0",
		16#516f# => X"ba050085",
		16#5170# => X"9dce0001",
		16#5171# => X"d7e117e8",
		16#5172# => X"d7e197f4",
		16#5173# => X"d7e1a7f8",
		16#5174# => X"84c40008",
		16#5175# => X"d7e14ffc",
		16#5176# => X"e1ce8000",
		16#5177# => X"a8440000",
		16#5178# => X"9c21ffe8",
		16#5179# => X"aa850000",
		16#517a# => X"aa430000",
		16#517b# => X"e5ae3000",
		16#517c# => X"10000006",
		16#517d# => X"84840004",
		16#517e# => X"e0c63000",
		16#517f# => X"e54e3000",
		16#5180# => X"13fffffe",
		16#5181# => X"9c840001",
		16#5182# => X"07fffdc7",
		16#5183# => X"a8720000",
		16#5184# => X"bdb00000",
		16#5185# => X"a90b0000",
		16#5186# => X"1000000c",
		16#5187# => X"9ccb0014",
		16#5188# => X"9ce00000",
		16#5189# => X"9c600000",
		16#518a# => X"9ce70001",
		16#518b# => X"d4061800",
		16#518c# => X"e4278000",
		16#518d# => X"13fffffd",
		16#518e# => X"9cc60004",
		16#518f# => X"9cc70005",
		16#5190# => X"b8c60002",
		16#5191# => X"e0c83000",
		16#5192# => X"85620010",
		16#5193# => X"a4b4001f",
		16#5194# => X"9d6b0005",
		16#5195# => X"9ce20014",
		16#5196# => X"b96b0002",
		16#5197# => X"bc050000",
		16#5198# => X"10000025",
		16#5199# => X"e1625800",
		16#519a# => X"9da00020",
		16#519b# => X"9c800000",
		16#519c# => X"e1ad2802",
		16#519d# => X"85870000",
		16#519e# => X"e18c2808",
		16#519f# => X"e0846004",
		16#51a0# => X"d4062000",
		16#51a1# => X"9cc60004",
		16#51a2# => X"84870000",
		16#51a3# => X"9ce70004",
		16#51a4# => X"e44b3800",
		16#51a5# => X"13fffff8",
		16#51a6# => X"e0846848",
		16#51a7# => X"bc040000",
		16#51a8# => X"10000003",
		16#51a9# => X"d4062000",
		16#51aa# => X"9dce0001",
		16#51ab# => X"84620004",
		16#51ac# => X"8492004c",
		16#51ad# => X"b8630002",
		16#51ae# => X"9dceffff",
		16#51af# => X"a9680000",
		16#51b0# => X"e0641800",
		16#51b1# => X"d4087010",
		16#51b2# => X"84830000",
		16#51b3# => X"d4022000",
		16#51b4# => X"d4031000",
		16#51b5# => X"9c210018",
		16#51b6# => X"8521fffc",
		16#51b7# => X"8441ffe8",
		16#51b8# => X"85c1ffec",
		16#51b9# => X"8601fff0",
		16#51ba# => X"8641fff4",
		16#51bb# => X"44004800",
		16#51bc# => X"8681fff8",
		16#51bd# => X"84670000",
		16#51be# => X"9ce70004",
		16#51bf# => X"d4061800",
		16#51c0# => X"e44b3800",
		16#51c1# => X"0fffffea",
		16#51c2# => X"9cc60004",
		16#51c3# => X"84670000",
		16#51c4# => X"9ce70004",
		16#51c5# => X"d4061800",
		16#51c6# => X"e44b3800",
		16#51c7# => X"13fffff6",
		16#51c8# => X"9cc60004",
		16#51c9# => X"03ffffe3",
		16#51ca# => X"84620004",
		16#51cb# => X"85630010",
		16#51cc# => X"84a40010",
		16#51cd# => X"e16b2802",
		16#51ce# => X"bc2b0000",
		16#51cf# => X"10000010",
		16#51d0# => X"15000000",
		16#51d1# => X"9ca50005",
		16#51d2# => X"9ce30014",
		16#51d3# => X"b8a50002",
		16#51d4# => X"e0632800",
		16#51d5# => X"e0842800",
		16#51d6# => X"9c63fffc",
		16#51d7# => X"9c84fffc",
		16#51d8# => X"84c30000",
		16#51d9# => X"84a40000",
		16#51da# => X"e4062800",
		16#51db# => X"0c000006",
		16#51dc# => X"e4871800",
		16#51dd# => X"13fffff9",
		16#51de# => X"15000000",
		16#51df# => X"44004800",
		16#51e0# => X"15000000",
		16#51e1# => X"e4662800",
		16#51e2# => X"13fffffd",
		16#51e3# => X"9d600001",
		16#51e4# => X"44004800",
		16#51e5# => X"9d60ffff",
		16#51e6# => X"d7e117ec",
		16#51e7# => X"a8440000",
		16#51e8# => X"d7e177f0",
		16#51e9# => X"d7e187f4",
		16#51ea# => X"d7e197f8",
		16#51eb# => X"d7e14ffc",
		16#51ec# => X"aa430000",
		16#51ed# => X"9c21ffec",
		16#51ee# => X"a8850000",
		16#51ef# => X"a8620000",
		16#51f0# => X"07ffffdb",
		16#51f1# => X"a9c50000",
		16#51f2# => X"bc2b0000",
		16#51f3# => X"0c00005a",
		16#51f4# => X"aa0b0000",
		16#51f5# => X"bd8b0000",
		16#51f6# => X"10000053",
		16#51f7# => X"9e000001",
		16#51f8# => X"9e000000",
		16#51f9# => X"a8720000",
		16#51fa# => X"07fffd4f",
		16#51fb# => X"84820004",
		16#51fc# => X"846e0010",
		16#51fd# => X"85820010",
		16#51fe# => X"9c630005",
		16#51ff# => X"9dec0005",
		16#5200# => X"b8630002",
		16#5201# => X"b9ef0002",
		16#5202# => X"9cee0014",
		16#5203# => X"d40b800c",
		16#5204# => X"e1ce1800",
		16#5205# => X"9cc20014",
		16#5206# => X"e1e27800",
		16#5207# => X"9c6b0014",
		16#5208# => X"9d000000",
		16#5209# => X"86a60000",
		16#520a# => X"86670000",
		16#520b# => X"a635ffff",
		16#520c# => X"a5b3ffff",
		16#520d# => X"bab50050",
		16#520e# => X"e1b16802",
		16#520f# => X"ba730050",
		16#5210# => X"e1ad4000",
		16#5211# => X"9ce70004",
		16#5212# => X"ba2d0090",
		16#5213# => X"e1159802",
		16#5214# => X"a5adffff",
		16#5215# => X"e1088800",
		16#5216# => X"9cc60004",
		16#5217# => X"ba280010",
		16#5218# => X"e44e3800",
		16#5219# => X"b9080090",
		16#521a# => X"e1b16804",
		16#521b# => X"d4036800",
		16#521c# => X"13ffffed",
		16#521d# => X"9c630004",
		16#521e# => X"a8430000",
		16#521f# => X"e4af3000",
		16#5220# => X"10000017",
		16#5221# => X"a8860000",
		16#5222# => X"84e60000",
		16#5223# => X"9cc60004",
		16#5224# => X"a4a7ffff",
		16#5225# => X"b8e70050",
		16#5226# => X"e0a82800",
		16#5227# => X"e44f3000",
		16#5228# => X"b9050090",
		16#5229# => X"a4a5ffff",
		16#522a# => X"e1083800",
		16#522b# => X"b8e80010",
		16#522c# => X"b9080090",
		16#522d# => X"e0a72804",
		16#522e# => X"d4032800",
		16#522f# => X"13fffff3",
		16#5230# => X"9c630004",
		16#5231# => X"ac64ffff",
		16#5232# => X"9c80fffc",
		16#5233# => X"e0637800",
		16#5234# => X"e0632003",
		16#5235# => X"9c630004",
		16#5236# => X"e0621800",
		16#5237# => X"9c63fffc",
		16#5238# => X"84430000",
		16#5239# => X"bc220000",
		16#523a# => X"10000007",
		16#523b# => X"15000000",
		16#523c# => X"9c63fffc",
		16#523d# => X"84430000",
		16#523e# => X"bc020000",
		16#523f# => X"13fffffd",
		16#5240# => X"9d8cffff",
		16#5241# => X"d40b6010",
		16#5242# => X"9c210014",
		16#5243# => X"8521fffc",
		16#5244# => X"8441ffec",
		16#5245# => X"85c1fff0",
		16#5246# => X"8601fff4",
		16#5247# => X"44004800",
		16#5248# => X"8641fff8",
		16#5249# => X"a8620000",
		16#524a# => X"a84e0000",
		16#524b# => X"03ffffae",
		16#524c# => X"a9c30000",
		16#524d# => X"a8720000",
		16#524e# => X"9c400001",
		16#524f# => X"07fffcfa",
		16#5250# => X"a88b0000",
		16#5251# => X"d40b8014",
		16#5252# => X"d40b1010",
		16#5253# => X"9c210014",
		16#5254# => X"8521fffc",
		16#5255# => X"8441ffec",
		16#5256# => X"85c1fff0",
		16#5257# => X"8601fff4",
		16#5258# => X"44004800",
		16#5259# => X"8641fff8",
		16#525a# => X"d7e117fc",
		16#525b# => X"18407ff0",
		16#525c# => X"9c21fffc",
		16#525d# => X"e0631003",
		16#525e# => X"1840fcc0",
		16#525f# => X"e0631000",
		16#5260# => X"bda30000",
		16#5261# => X"10000007",
		16#5262# => X"9c800000",
		16#5263# => X"9c210004",
		16#5264# => X"a9630000",
		16#5265# => X"a9840000",
		16#5266# => X"44004800",
		16#5267# => X"8441fffc",
		16#5268# => X"e0601802",
		16#5269# => X"b8630094",
		16#526a# => X"bd430013",
		16#526b# => X"0c00000e",
		16#526c# => X"9ca3ffec",
		16#526d# => X"9c800001",
		16#526e# => X"bd45001e",
		16#526f# => X"13fffff4",
		16#5270# => X"9c600000",
		16#5271# => X"9cc0001f",
		16#5272# => X"9c210004",
		16#5273# => X"e0a62802",
		16#5274# => X"a9630000",
		16#5275# => X"e0842808",
		16#5276# => X"8441fffc",
		16#5277# => X"44004800",
		16#5278# => X"a9840000",
		16#5279# => X"18a00008",
		16#527a# => X"9c800000",
		16#527b# => X"e0651888",
		16#527c# => X"9c210004",
		16#527d# => X"a9840000",
		16#527e# => X"a9630000",
		16#527f# => X"44004800",
		16#5280# => X"8441fffc",
		16#5281# => X"d7e197f4",
		16#5282# => X"86430010",
		16#5283# => X"d7e117e8",
		16#5284# => X"9e520005",
		16#5285# => X"d7e177ec",
		16#5286# => X"ba520002",
		16#5287# => X"d7e187f0",
		16#5288# => X"d7e1a7f8",
		16#5289# => X"e2439000",
		16#528a# => X"d7e14ffc",
		16#528b# => X"9c52fffc",
		16#528c# => X"9c21ffe8",
		16#528d# => X"85c20000",
		16#528e# => X"9e030014",
		16#528f# => X"a86e0000",
		16#5290# => X"07fffd82",
		16#5291# => X"aa840000",
		16#5292# => X"9c600020",
		16#5293# => X"bd4b000a",
		16#5294# => X"e0635802",
		16#5295# => X"10000019",
		16#5296# => X"d4141800",
		16#5297# => X"9ca0000b",
		16#5298# => X"18c03ff0",
		16#5299# => X"e0a55802",
		16#529a# => X"9c800000",
		16#529b# => X"e06e2848",
		16#529c# => X"e4701000",
		16#529d# => X"10000004",
		16#529e# => X"e0633004",
		16#529f# => X"8482fffc",
		16#52a0# => X"e0842848",
		16#52a1# => X"9d6b0015",
		16#52a2# => X"e1ce5808",
		16#52a3# => X"e1c47004",
		16#52a4# => X"9c210018",
		16#52a5# => X"a98e0000",
		16#52a6# => X"8521fffc",
		16#52a7# => X"a9630000",
		16#52a8# => X"8441ffe8",
		16#52a9# => X"85c1ffec",
		16#52aa# => X"8601fff0",
		16#52ab# => X"8641fff4",
		16#52ac# => X"44004800",
		16#52ad# => X"8681fff8",
		16#52ae# => X"e4701000",
		16#52af# => X"10000004",
		16#52b0# => X"9c800000",
		16#52b1# => X"9c52fff8",
		16#52b2# => X"84820000",
		16#52b3# => X"9d6bfff5",
		16#52b4# => X"bc0b0000",
		16#52b5# => X"10000010",
		16#52b6# => X"19003ff0",
		16#52b7# => X"9cc00020",
		16#52b8# => X"e06e5808",
		16#52b9# => X"e0c65802",
		16#52ba# => X"e0e43048",
		16#52bb# => X"e0634004",
		16#52bc# => X"9ca00000",
		16#52bd# => X"e4a28000",
		16#52be# => X"10000004",
		16#52bf# => X"e0633804",
		16#52c0# => X"84a2fffc",
		16#52c1# => X"e0a53048",
		16#52c2# => X"e1c45808",
		16#52c3# => X"03ffffe1",
		16#52c4# => X"e1c57004",
		16#52c5# => X"18403ff0",
		16#52c6# => X"e06e1004",
		16#52c7# => X"03ffffdd",
		16#52c8# => X"a9c40000",
		16#52c9# => X"d7e117e4",
		16#52ca# => X"d7e177e8",
		16#52cb# => X"d7e187ec",
		16#52cc# => X"d7e197f0",
		16#52cd# => X"d7e1a7f4",
		16#52ce# => X"d7e1b7f8",
		16#52cf# => X"aa040000",
		16#52d0# => X"d7e14ffc",
		16#52d1# => X"9c800001",
		16#52d2# => X"9c21ffdc",
		16#52d3# => X"aac60000",
		16#52d4# => X"aa870000",
		16#52d5# => X"07fffc74",
		16#52d6# => X"aa450000",
		16#52d7# => X"18607fff",
		16#52d8# => X"a84b0000",
		16#52d9# => X"a863ffff",
		16#52da# => X"e1d01803",
		16#52db# => X"1860000f",
		16#52dc# => X"b9ce0054",
		16#52dd# => X"a863ffff",
		16#52de# => X"e2101803",
		16#52df# => X"bc0e0000",
		16#52e0# => X"10000005",
		16#52e1# => X"d4018000",
		16#52e2# => X"18600010",
		16#52e3# => X"e2101804",
		16#52e4# => X"d4018000",
		16#52e5# => X"bc120000",
		16#52e6# => X"1000001a",
		16#52e7# => X"a8610000",
		16#52e8# => X"9c610004",
		16#52e9# => X"07fffd54",
		16#52ea# => X"d4019004",
		16#52eb# => X"bc0b0000",
		16#52ec# => X"0c000030",
		16#52ed# => X"9c800020",
		16#52ee# => X"84810004",
		16#52ef# => X"84610000",
		16#52f0# => X"d4022014",
		16#52f1# => X"d4021818",
		16#52f2# => X"bc030000",
		16#52f3# => X"10000003",
		16#52f4# => X"9e000001",
		16#52f5# => X"9e000002",
		16#52f6# => X"bc0e0000",
		16#52f7# => X"10000011",
		16#52f8# => X"d4028010",
		16#52f9# => X"9dcefbcd",
		16#52fa# => X"9c600035",
		16#52fb# => X"e1ce5800",
		16#52fc# => X"e1635802",
		16#52fd# => X"d4167000",
		16#52fe# => X"00000014",
		16#52ff# => X"d4145800",
		16#5300# => X"07fffd3d",
		16#5301# => X"9e000001",
		16#5302# => X"84610000",
		16#5303# => X"d4028010",
		16#5304# => X"d4021814",
		16#5305# => X"bc0e0000",
		16#5306# => X"0ffffff3",
		16#5307# => X"9d6b0020",
		16#5308# => X"9c700004",
		16#5309# => X"9d6bfbce",
		16#530a# => X"b8630002",
		16#530b# => X"ba100005",
		16#530c# => X"d4165800",
		16#530d# => X"e0621800",
		16#530e# => X"07fffd04",
		16#530f# => X"84630000",
		16#5310# => X"e1705802",
		16#5311# => X"d4145800",
		16#5312# => X"9c210024",
		16#5313# => X"a9620000",
		16#5314# => X"8521fffc",
		16#5315# => X"8441ffe4",
		16#5316# => X"85c1ffe8",
		16#5317# => X"8601ffec",
		16#5318# => X"8641fff0",
		16#5319# => X"8681fff4",
		16#531a# => X"44004800",
		16#531b# => X"86c1fff8",
		16#531c# => X"84610000",
		16#531d# => X"e0845802",
		16#531e# => X"84a10004",
		16#531f# => X"e0832008",
		16#5320# => X"e0635848",
		16#5321# => X"e0842804",
		16#5322# => X"d4011800",
		16#5323# => X"03ffffce",
		16#5324# => X"d4022014",
		16#5325# => X"d7e14ffc",
		16#5326# => X"d7e117e4",
		16#5327# => X"d7e177e8",
		16#5328# => X"d7e187ec",
		16#5329# => X"d7e197f0",
		16#532a# => X"d7e1a7f4",
		16#532b# => X"d7e1b7f8",
		16#532c# => X"9c21ffdc",
		16#532d# => X"aa440000",
		16#532e# => X"9c810004",
		16#532f# => X"07ffff52",
		16#5330# => X"aa830000",
		16#5331# => X"a8720000",
		16#5332# => X"a8810000",
		16#5333# => X"a9cb0000",
		16#5334# => X"07ffff4d",
		16#5335# => X"aa0c0000",
		16#5336# => X"84740010",
		16#5337# => X"84920010",
		16#5338# => X"84a10004",
		16#5339# => X"e0832002",
		16#533a# => X"84610000",
		16#533b# => X"b8840005",
		16#533c# => X"e0651802",
		16#533d# => X"a84b0000",
		16#533e# => X"e0632000",
		16#533f# => X"aace0000",
		16#5340# => X"a8ec0000",
		16#5341# => X"bda30000",
		16#5342# => X"10000016",
		16#5343# => X"a8a20000",
		16#5344# => X"b9c30014",
		16#5345# => X"e1ceb000",
		16#5346# => X"a86e0000",
		16#5347# => X"a8a20000",
		16#5348# => X"a8900000",
		16#5349# => X"07ffdac3",
		16#534a# => X"a8c70000",
		16#534b# => X"9c210024",
		16#534c# => X"a84b0000",
		16#534d# => X"a86c0000",
		16#534e# => X"8521fffc",
		16#534f# => X"e1620004",
		16#5350# => X"e1830004",
		16#5351# => X"85c1ffe8",
		16#5352# => X"8441ffe4",
		16#5353# => X"8601ffec",
		16#5354# => X"8641fff0",
		16#5355# => X"8681fff4",
		16#5356# => X"44004800",
		16#5357# => X"86c1fff8",
		16#5358# => X"b8430014",
		16#5359# => X"03ffffed",
		16#535a# => X"e0451002",
		16#535b# => X"d7e117f8",
		16#535c# => X"d7e14ffc",
		16#535d# => X"a8430000",
		16#535e# => X"bd430017",
		16#535f# => X"0c000017",
		16#5360# => X"9c21fff8",
		16#5361# => X"19603ff0",
		16#5362# => X"9d800000",
		16#5363# => X"18e00001",
		16#5364# => X"a86b0000",
		16#5365# => X"a8e78afc",
		16#5366# => X"a88c0000",
		16#5367# => X"84a70000",
		16#5368# => X"84c70004",
		16#5369# => X"07ffd9a0",
		16#536a# => X"9c42ffff",
		16#536b# => X"bc220000",
		16#536c# => X"13fffff8",
		16#536d# => X"18e00001",
		16#536e# => X"9c210008",
		16#536f# => X"a84b0000",
		16#5370# => X"a86c0000",
		16#5371# => X"8521fffc",
		16#5372# => X"e1620004",
		16#5373# => X"e1830004",
		16#5374# => X"44004800",
		16#5375# => X"8441fff8",
		16#5376# => X"b8430003",
		16#5377# => X"18600001",
		16#5378# => X"9c210008",
		16#5379# => X"a8638b04",
		16#537a# => X"8521fffc",
		16#537b# => X"e0421800",
		16#537c# => X"85820004",
		16#537d# => X"85620000",
		16#537e# => X"a86c0000",
		16#537f# => X"a84b0000",
		16#5380# => X"e1620004",
		16#5381# => X"e1830004",
		16#5382# => X"44004800",
		16#5383# => X"8441fff8",
		16#5384# => X"9c84ffff",
		16#5385# => X"84e50010",
		16#5386# => X"b9040085",
		16#5387# => X"9ce70005",
		16#5388# => X"d7e117fc",
		16#5389# => X"9d080001",
		16#538a# => X"b8e70002",
		16#538b# => X"b9080002",
		16#538c# => X"9c850014",
		16#538d# => X"e0e53800",
		16#538e# => X"9c21fffc",
		16#538f# => X"e4643800",
		16#5390# => X"1000000f",
		16#5391# => X"e1034000",
		16#5392# => X"a8c30000",
		16#5393# => X"85640000",
		16#5394# => X"9c840004",
		16#5395# => X"d4065800",
		16#5396# => X"e4472000",
		16#5397# => X"13fffffc",
		16#5398# => X"9cc60004",
		16#5399# => X"e0872802",
		16#539a# => X"9c40fffc",
		16#539b# => X"9c84ffeb",
		16#539c# => X"e0841003",
		16#539d# => X"9c840004",
		16#539e# => X"e0632000",
		16#539f# => X"e4a81800",
		16#53a0# => X"10000008",
		16#53a1# => X"15000000",
		16#53a2# => X"9c400000",
		16#53a3# => X"d4031000",
		16#53a4# => X"9c630004",
		16#53a5# => X"e4481800",
		16#53a6# => X"13fffffd",
		16#53a7# => X"15000000",
		16#53a8# => X"9c210004",
		16#53a9# => X"44004800",
		16#53aa# => X"8441fffc",
		16#53ab# => X"b8a40085",
		16#53ac# => X"84c30010",
		16#53ad# => X"e5662800",
		16#53ae# => X"10000019",
		16#53af# => X"e5462800",
		16#53b0# => X"a8a60000",
		16#53b1# => X"9ca50005",
		16#53b2# => X"9c830014",
		16#53b3# => X"b8a50002",
		16#53b4# => X"e0632800",
		16#53b5# => X"e4641800",
		16#53b6# => X"1000000f",
		16#53b7# => X"9d600000",
		16#53b8# => X"9c63fffc",
		16#53b9# => X"84a30000",
		16#53ba# => X"bc250000",
		16#53bb# => X"1000000a",
		16#53bc# => X"9d600001",
		16#53bd# => X"e4841800",
		16#53be# => X"0c000018",
		16#53bf# => X"9c63fffc",
		16#53c0# => X"84a30000",
		16#53c1# => X"bc250000",
		16#53c2# => X"0ffffffc",
		16#53c3# => X"e4841800",
		16#53c4# => X"9d600001",
		16#53c5# => X"44004800",
		16#53c6# => X"15000000",
		16#53c7# => X"0fffffea",
		16#53c8# => X"a484001f",
		16#53c9# => X"bc240000",
		16#53ca# => X"0fffffe7",
		16#53cb# => X"9cc50005",
		16#53cc# => X"b8c60002",
		16#53cd# => X"e0c33000",
		16#53ce# => X"84c60000",
		16#53cf# => X"e0e62048",
		16#53d0# => X"e0872008",
		16#53d1# => X"e4243000",
		16#53d2# => X"0fffffdf",
		16#53d3# => X"9d600001",
		16#53d4# => X"44004800",
		16#53d5# => X"15000000",
		16#53d6# => X"44004800",
		16#53d7# => X"9d600000",
		16#53d8# => X"d7e187dc",
		16#53d9# => X"d7e197e0",
		16#53da# => X"d7e1c7ec",
		16#53db# => X"d7e14ffc",
		16#53dc# => X"d7e117d4",
		16#53dd# => X"d7e177d8",
		16#53de# => X"d7e1a7e4",
		16#53df# => X"d7e1b7e8",
		16#53e0# => X"d7e1d7f0",
		16#53e1# => X"d7e1e7f4",
		16#53e2# => X"d7e1f7f8",
		16#53e3# => X"aa040000",
		16#53e4# => X"9c21ffd4",
		16#53e5# => X"ab030000",
		16#53e6# => X"bc240000",
		16#53e7# => X"0c00010f",
		16#53e8# => X"aa450000",
		16#53e9# => X"9c50fff8",
		16#53ea# => X"07ffdff0",
		16#53eb# => X"9dd2000b",
		16#53ec# => X"bcae0016",
		16#53ed# => X"0c000065",
		16#53ee# => X"84c20004",
		16#53ef# => X"9c600010",
		16#53f0# => X"9c800000",
		16#53f1# => X"a9c30000",
		16#53f2# => X"e48e9000",
		16#53f3# => X"10000003",
		16#53f4# => X"9ca00001",
		16#53f5# => X"9ca00000",
		16#53f6# => X"a4a500ff",
		16#53f7# => X"bc250000",
		16#53f8# => X"1000010c",
		16#53f9# => X"bc040000",
		16#53fa# => X"0c00010a",
		16#53fb# => X"9ca0fffc",
		16#53fc# => X"e2862803",
		16#53fd# => X"e5741800",
		16#53fe# => X"10000059",
		16#53ff# => X"aad40000",
		16#5400# => X"1b800001",
		16#5401# => X"e0e2a000",
		16#5402# => X"ab9cb20c",
		16#5403# => X"84bc0008",
		16#5404# => X"e4053800",
		16#5405# => X"10000103",
		16#5406# => X"9d80fffe",
		16#5407# => X"85070004",
		16#5408# => X"e1686003",
		16#5409# => X"e1675800",
		16#540a# => X"856b0004",
		16#540b# => X"a56b0001",
		16#540c# => X"bc0b0000",
		16#540d# => X"10000066",
		16#540e# => X"9d60fffc",
		16#540f# => X"a8e40000",
		16#5410# => X"a4c60001",
		16#5411# => X"bc260000",
		16#5412# => X"1000007a",
		16#5413# => X"9d60fffc",
		16#5414# => X"87420000",
		16#5415# => X"e342d002",
		16#5416# => X"bc070000",
		16#5417# => X"87da0004",
		16#5418# => X"100000ad",
		16#5419# => X"e3de5803",
		16#541a# => X"e4272800",
		16#541b# => X"0c00010f",
		16#541c# => X"9cae0010",
		16#541d# => X"e3dea000",
		16#541e# => X"e2c4f000",
		16#541f# => X"e543b000",
		16#5420# => X"100000a7",
		16#5421# => X"e543f000",
		16#5422# => X"8447000c",
		16#5423# => X"84670008",
		16#5424# => X"9cb4fffc",
		16#5425# => X"d403100c",
		16#5426# => X"d4021808",
		16#5427# => X"845a000c",
		16#5428# => X"847a0008",
		16#5429# => X"9e5a0008",
		16#542a# => X"d403100c",
		16#542b# => X"bc450024",
		16#542c# => X"1000013f",
		16#542d# => X"d4021808",
		16#542e# => X"bca50013",
		16#542f# => X"10000018",
		16#5430# => X"a8520000",
		16#5431# => X"84700000",
		16#5432# => X"9c5a0010",
		16#5433# => X"d4121800",
		16#5434# => X"bca5001b",
		16#5435# => X"84700004",
		16#5436# => X"9e100008",
		16#5437# => X"10000010",
		16#5438# => X"d41a180c",
		16#5439# => X"84700000",
		16#543a# => X"bc250024",
		16#543b# => X"d4021800",
		16#543c# => X"9c5a0018",
		16#543d# => X"84700004",
		16#543e# => X"9e100008",
		16#543f# => X"10000008",
		16#5440# => X"d41a1814",
		16#5441# => X"84700000",
		16#5442# => X"d4021800",
		16#5443# => X"9c5a0020",
		16#5444# => X"84700004",
		16#5445# => X"9e100008",
		16#5446# => X"d41a181c",
		16#5447# => X"84700000",
		16#5448# => X"9e100004",
		16#5449# => X"d4021800",
		16#544a# => X"9c620004",
		16#544b# => X"84500000",
		16#544c# => X"d4031000",
		16#544d# => X"a85a0000",
		16#544e# => X"84900004",
		16#544f# => X"d4032004",
		16#5450# => X"00000008",
		16#5451# => X"84da0004",
		16#5452# => X"9c60fff8",
		16#5453# => X"e1ce1803",
		16#5454# => X"a86e0000",
		16#5455# => X"03ffff9d",
		16#5456# => X"b88e005f",
		16#5457# => X"9e420008",
		16#5458# => X"e0767002",
		16#5459# => X"bca3000f",
		16#545a# => X"0c000024",
		16#545b# => X"e0827000",
		16#545c# => X"a4c60001",
		16#545d# => X"e062b000",
		16#545e# => X"e2c6b004",
		16#545f# => X"d402b004",
		16#5460# => X"84430004",
		16#5461# => X"a8420001",
		16#5462# => X"d4031004",
		16#5463# => X"07ffdf79",
		16#5464# => X"a8780000",
		16#5465# => X"9c21002c",
		16#5466# => X"a9720000",
		16#5467# => X"8521fffc",
		16#5468# => X"8441ffd4",
		16#5469# => X"85c1ffd8",
		16#546a# => X"8601ffdc",
		16#546b# => X"8641ffe0",
		16#546c# => X"8681ffe4",
		16#546d# => X"86c1ffe8",
		16#546e# => X"8701ffec",
		16#546f# => X"8741fff0",
		16#5470# => X"8781fff4",
		16#5471# => X"44004800",
		16#5472# => X"87c1fff8",
		16#5473# => X"e0885803",
		16#5474# => X"e2c4a000",
		16#5475# => X"e5a3b000",
		16#5476# => X"0fffff9a",
		16#5477# => X"15000000",
		16#5478# => X"8467000c",
		16#5479# => X"84870008",
		16#547a# => X"9e420008",
		16#547b# => X"d404180c",
		16#547c# => X"03ffffdc",
		16#547d# => X"d4032008",
		16#547e# => X"a4c60001",
		16#547f# => X"e1c67004",
		16#5480# => X"a8a30001",
		16#5481# => X"d4027004",
		16#5482# => X"d4042804",
		16#5483# => X"e0441800",
		16#5484# => X"a8780000",
		16#5485# => X"84a20004",
		16#5486# => X"9c840008",
		16#5487# => X"a8a50001",
		16#5488# => X"07fff627",
		16#5489# => X"d4022804",
		16#548a# => X"03ffffd9",
		16#548b# => X"15000000",
		16#548c# => X"a8920000",
		16#548d# => X"07ffdcfd",
		16#548e# => X"a8780000",
		16#548f# => X"bc2b0000",
		16#5490# => X"0fffffd3",
		16#5491# => X"aa4b0000",
		16#5492# => X"84c20004",
		16#5493# => X"9d80fffe",
		16#5494# => X"9c6bfff8",
		16#5495# => X"e0866003",
		16#5496# => X"e0822000",
		16#5497# => X"e4232000",
		16#5498# => X"0c0000cd",
		16#5499# => X"9cb4fffc",
		16#549a# => X"bc450024",
		16#549b# => X"1000008a",
		16#549c# => X"a8500000",
		16#549d# => X"bca50013",
		16#549e# => X"10000018",
		16#549f# => X"a86b0000",
		16#54a0# => X"84500000",
		16#54a1# => X"9c6b0008",
		16#54a2# => X"d40b1000",
		16#54a3# => X"bca5001b",
		16#54a4# => X"84900004",
		16#54a5# => X"9c500008",
		16#54a6# => X"10000010",
		16#54a7# => X"d40b2004",
		16#54a8# => X"84420000",
		16#54a9# => X"bc250024",
		16#54aa# => X"d4031000",
		16#54ab# => X"9c500010",
		16#54ac# => X"8490000c",
		16#54ad# => X"9c6b0010",
		16#54ae# => X"10000008",
		16#54af# => X"d40b200c",
		16#54b0# => X"84820000",
		16#54b1# => X"9c500018",
		16#54b2# => X"d4032000",
		16#54b3# => X"9c6b0018",
		16#54b4# => X"84900014",
		16#54b5# => X"d40b2014",
		16#54b6# => X"84820000",
		16#54b7# => X"9c420004",
		16#54b8# => X"d4032000",
		16#54b9# => X"9c630004",
		16#54ba# => X"84820000",
		16#54bb# => X"d4032000",
		16#54bc# => X"84420004",
		16#54bd# => X"d4031004",
		16#54be# => X"a8780000",
		16#54bf# => X"07fff5f0",
		16#54c0# => X"a8900000",
		16#54c1# => X"07ffdf1b",
		16#54c2# => X"a8780000",
		16#54c3# => X"03ffffa3",
		16#54c4# => X"9c21002c",
		16#54c5# => X"e3dea000",
		16#54c6# => X"e543f000",
		16#54c7# => X"13ffffc6",
		16#54c8# => X"a8920000",
		16#54c9# => X"845a000c",
		16#54ca# => X"847a0008",
		16#54cb# => X"9cb4fffc",
		16#54cc# => X"d403100c",
		16#54cd# => X"d4021808",
		16#54ce# => X"bc450024",
		16#54cf# => X"1000004f",
		16#54d0# => X"9e5a0008",
		16#54d1# => X"bca50013",
		16#54d2# => X"10000018",
		16#54d3# => X"a8520000",
		16#54d4# => X"84700000",
		16#54d5# => X"9c5a0010",
		16#54d6# => X"d4121800",
		16#54d7# => X"bca5001b",
		16#54d8# => X"84700004",
		16#54d9# => X"9e100008",
		16#54da# => X"10000010",
		16#54db# => X"d41a180c",
		16#54dc# => X"84700000",
		16#54dd# => X"bc250024",
		16#54de# => X"d4021800",
		16#54df# => X"9c5a0018",
		16#54e0# => X"84700004",
		16#54e1# => X"9e100008",
		16#54e2# => X"10000008",
		16#54e3# => X"d41a1814",
		16#54e4# => X"84700000",
		16#54e5# => X"d4021800",
		16#54e6# => X"9c5a0020",
		16#54e7# => X"84700004",
		16#54e8# => X"9e100008",
		16#54e9# => X"d41a181c",
		16#54ea# => X"84700000",
		16#54eb# => X"9e100004",
		16#54ec# => X"d4021800",
		16#54ed# => X"9c620004",
		16#54ee# => X"84500000",
		16#54ef# => X"aade0000",
		16#54f0# => X"d4031000",
		16#54f1# => X"a85a0000",
		16#54f2# => X"84900004",
		16#54f3# => X"d4032004",
		16#54f4# => X"03ffff64",
		16#54f5# => X"84da0004",
		16#54f6# => X"9c21002c",
		16#54f7# => X"a8850000",
		16#54f8# => X"8521fffc",
		16#54f9# => X"8441ffd4",
		16#54fa# => X"85c1ffd8",
		16#54fb# => X"8601ffdc",
		16#54fc# => X"8641ffe0",
		16#54fd# => X"8681ffe4",
		16#54fe# => X"86c1ffe8",
		16#54ff# => X"8701ffec",
		16#5500# => X"8741fff0",
		16#5501# => X"8781fff4",
		16#5502# => X"03ffdc88",
		16#5503# => X"87c1fff8",
		16#5504# => X"9c40000c",
		16#5505# => X"9e400000",
		16#5506# => X"03ffff5f",
		16#5507# => X"d4181000",
		16#5508# => X"9ce0fffc",
		16#5509# => X"84850004",
		16#550a# => X"9d6e0010",
		16#550b# => X"e0843803",
		16#550c# => X"e104a000",
		16#550d# => X"e5885800",
		16#550e# => X"13ffff02",
		16#550f# => X"a8e50000",
		16#5510# => X"e0a87002",
		16#5511# => X"e0827000",
		16#5512# => X"a8a50001",
		16#5513# => X"d41c2008",
		16#5514# => X"d4042804",
		16#5515# => X"a8780000",
		16#5516# => X"84820004",
		16#5517# => X"aa500000",
		16#5518# => X"a4840001",
		16#5519# => X"e1ce2004",
		16#551a# => X"07ffdec2",
		16#551b# => X"d4027004",
		16#551c# => X"03ffff4a",
		16#551d# => X"9c21002c",
		16#551e# => X"a8720000",
		16#551f# => X"a8900000",
		16#5520# => X"07fff97a",
		16#5521# => X"aade0000",
		16#5522# => X"84da0004",
		16#5523# => X"03ffff35",
		16#5524# => X"a85a0000",
		16#5525# => X"a86b0000",
		16#5526# => X"07fff974",
		16#5527# => X"a8900000",
		16#5528# => X"03ffff97",
		16#5529# => X"a8780000",
		16#552a# => X"e3dea000",
		16#552b# => X"e2c4f000",
		16#552c# => X"e5962800",
		16#552d# => X"13ffff9a",
		16#552e# => X"e543f000",
		16#552f# => X"845a000c",
		16#5530# => X"847a0008",
		16#5531# => X"e0b45800",
		16#5532# => X"d403100c",
		16#5533# => X"d4021808",
		16#5534# => X"bc450024",
		16#5535# => X"1000003c",
		16#5536# => X"9e5a0008",
		16#5537# => X"bca50013",
		16#5538# => X"10000018",
		16#5539# => X"a8520000",
		16#553a# => X"84700000",
		16#553b# => X"9c5a0010",
		16#553c# => X"d4121800",
		16#553d# => X"bca5001b",
		16#553e# => X"84700004",
		16#553f# => X"9e100008",
		16#5540# => X"10000010",
		16#5541# => X"d41a180c",
		16#5542# => X"84700000",
		16#5543# => X"bc250024",
		16#5544# => X"d4021800",
		16#5545# => X"9c5a0018",
		16#5546# => X"84700004",
		16#5547# => X"9e100008",
		16#5548# => X"10000008",
		16#5549# => X"d41a1814",
		16#554a# => X"84700000",
		16#554b# => X"d4021800",
		16#554c# => X"9c5a0020",
		16#554d# => X"84700004",
		16#554e# => X"9e100008",
		16#554f# => X"d41a181c",
		16#5550# => X"84700000",
		16#5551# => X"9e100004",
		16#5552# => X"d4021800",
		16#5553# => X"9c420004",
		16#5554# => X"84700000",
		16#5555# => X"d4021800",
		16#5556# => X"84700004",
		16#5557# => X"d4021804",
		16#5558# => X"e0967002",
		16#5559# => X"e05a7000",
		16#555a# => X"a8840001",
		16#555b# => X"d41c1008",
		16#555c# => X"d4022004",
		16#555d# => X"a8780000",
		16#555e# => X"845a0004",
		16#555f# => X"a4420001",
		16#5560# => X"e1ce1004",
		16#5561# => X"07ffde7b",
		16#5562# => X"d41a7004",
		16#5563# => X"03ffff03",
		16#5564# => X"9c21002c",
		16#5565# => X"86c30004",
		16#5566# => X"9c60fffc",
		16#5567# => X"9e420008",
		16#5568# => X"e2d61803",
		16#5569# => X"03fffeef",
		16#556a# => X"e2d6a000",
		16#556b# => X"a8720000",
		16#556c# => X"a8900000",
		16#556d# => X"07fff92d",
		16#556e# => X"a85a0000",
		16#556f# => X"03fffee9",
		16#5570# => X"84da0004",
		16#5571# => X"a8720000",
		16#5572# => X"07fff928",
		16#5573# => X"a8900000",
		16#5574# => X"03ffffe5",
		16#5575# => X"e0967002",
		16#5576# => X"d7e117f4",
		16#5577# => X"d7e177f8",
		16#5578# => X"d7e14ffc",
		16#5579# => X"a8440000",
		16#557a# => X"84840000",
		16#557b# => X"9c21fff4",
		16#557c# => X"bc040000",
		16#557d# => X"10000004",
		16#557e# => X"a9c30000",
		16#557f# => X"07fffff7",
		16#5580# => X"15000000",
		16#5581# => X"9c21000c",
		16#5582# => X"a86e0000",
		16#5583# => X"a8820000",
		16#5584# => X"8521fffc",
		16#5585# => X"8441fff4",
		16#5586# => X"03fff529",
		16#5587# => X"85c1fff8",
		16#5588# => X"d7e117ec",
		16#5589# => X"18400001",
		16#558a# => X"d7e177f0",
		16#558b# => X"a842ade4",
		16#558c# => X"d7e14ffc",
		16#558d# => X"d7e187f4",
		16#558e# => X"d7e197f8",
		16#558f# => X"84420000",
		16#5590# => X"9c21ffec",
		16#5591# => X"e4031000",
		16#5592# => X"1000003a",
		16#5593# => X"a9c30000",
		16#5594# => X"8483004c",
		16#5595# => X"bc040000",
		16#5596# => X"10000017",
		16#5597# => X"9c400000",
		16#5598# => X"aa020000",
		16#5599# => X"b8420002",
		16#559a# => X"e0441000",
		16#559b# => X"84a20000",
		16#559c# => X"bc050000",
		16#559d# => X"1000000a",
		16#559e# => X"15000000",
		16#559f# => X"a8850000",
		16#55a0# => X"a86e0000",
		16#55a1# => X"07fff50e",
		16#55a2# => X"84450000",
		16#55a3# => X"bc220000",
		16#55a4# => X"13fffffb",
		16#55a5# => X"a8a20000",
		16#55a6# => X"848e004c",
		16#55a7# => X"9e100001",
		16#55a8# => X"bc100020",
		16#55a9# => X"0ffffff0",
		16#55aa# => X"a8500000",
		16#55ab# => X"07fff504",
		16#55ac# => X"a86e0000",
		16#55ad# => X"848e0040",
		16#55ae# => X"bc040000",
		16#55af# => X"10000004",
		16#55b0# => X"15000000",
		16#55b1# => X"07fff4fe",
		16#55b2# => X"a86e0000",
		16#55b3# => X"844e0148",
		16#55b4# => X"bc020000",
		16#55b5# => X"1000000d",
		16#55b6# => X"15000000",
		16#55b7# => X"9e4e014c",
		16#55b8# => X"e4029000",
		16#55b9# => X"10000009",
		16#55ba# => X"15000000",
		16#55bb# => X"a8820000",
		16#55bc# => X"a86e0000",
		16#55bd# => X"07fff4f2",
		16#55be# => X"86020000",
		16#55bf# => X"e4328000",
		16#55c0# => X"13fffffb",
		16#55c1# => X"a8500000",
		16#55c2# => X"848e0054",
		16#55c3# => X"bc040000",
		16#55c4# => X"10000004",
		16#55c5# => X"15000000",
		16#55c6# => X"07fff4e9",
		16#55c7# => X"a86e0000",
		16#55c8# => X"844e0038",
		16#55c9# => X"bc020000",
		16#55ca# => X"0c000009",
		16#55cb# => X"15000000",
		16#55cc# => X"9c210014",
		16#55cd# => X"8521fffc",
		16#55ce# => X"8441ffec",
		16#55cf# => X"85c1fff0",
		16#55d0# => X"8601fff4",
		16#55d1# => X"44004800",
		16#55d2# => X"8641fff8",
		16#55d3# => X"844e003c",
		16#55d4# => X"48001000",
		16#55d5# => X"a86e0000",
		16#55d6# => X"848e02e0",
		16#55d7# => X"bc040000",
		16#55d8# => X"13fffff4",
		16#55d9# => X"15000000",
		16#55da# => X"9c210014",
		16#55db# => X"a86e0000",
		16#55dc# => X"8521fffc",
		16#55dd# => X"8441ffec",
		16#55de# => X"85c1fff0",
		16#55df# => X"8601fff4",
		16#55e0# => X"03ffff96",
		16#55e1# => X"8641fff8",
		16#55e2# => X"d7e197f8",
		16#55e3# => X"d7e14ffc",
		16#55e4# => X"d7e117ec",
		16#55e5# => X"d7e177f0",
		16#55e6# => X"d7e187f4",
		16#55e7# => X"aa430000",
		16#55e8# => X"bc230000",
		16#55e9# => X"0c000029",
		16#55ea# => X"9c21ffec",
		16#55eb# => X"86120148",
		16#55ec# => X"bc100000",
		16#55ed# => X"10000013",
		16#55ee# => X"15000000",
		16#55ef# => X"84500004",
		16#55f0# => X"9dc2ffff",
		16#55f1# => X"bd8e0000",
		16#55f2# => X"1000000a",
		16#55f3# => X"9c420001",
		16#55f4# => X"b8420002",
		16#55f5# => X"e0501000",
		16#55f6# => X"84820000",
		16#55f7# => X"48002000",
		16#55f8# => X"9dceffff",
		16#55f9# => X"bd6e0000",
		16#55fa# => X"13fffffc",
		16#55fb# => X"9c42fffc",
		16#55fc# => X"86100000",
		16#55fd# => X"bc300000",
		16#55fe# => X"13fffff1",
		16#55ff# => X"15000000",
		16#5600# => X"8452003c",
		16#5601# => X"bc020000",
		16#5602# => X"10000009",
		16#5603# => X"a8720000",
		16#5604# => X"9c210014",
		16#5605# => X"8521fffc",
		16#5606# => X"85c1fff0",
		16#5607# => X"8601fff4",
		16#5608# => X"8641fff8",
		16#5609# => X"44001000",
		16#560a# => X"8441ffec",
		16#560b# => X"9c210014",
		16#560c# => X"8521fffc",
		16#560d# => X"8441ffec",
		16#560e# => X"85c1fff0",
		16#560f# => X"8601fff4",
		16#5610# => X"44004800",
		16#5611# => X"8641fff8",
		16#5612# => X"18400001",
		16#5613# => X"a842ade4",
		16#5614# => X"03ffffd7",
		16#5615# => X"86420000",
		16#5616# => X"d7e117fc",
		16#5617# => X"e0a41804",
		16#5618# => X"9c21fffc",
		16#5619# => X"bc050000",
		16#561a# => X"10000041",
		16#561b# => X"9d600002",
		16#561c# => X"e0a02002",
		16#561d# => X"e0852004",
		16#561e# => X"ac84ffff",
		16#561f# => X"b884005f",
		16#5620# => X"bc040000",
		16#5621# => X"0c00003d",
		16#5622# => X"18408000",
		16#5623# => X"18407ff0",
		16#5624# => X"e0c31000",
		16#5625# => X"18407fdf",
		16#5626# => X"a842ffff",
		16#5627# => X"e4a61000",
		16#5628# => X"10000003",
		16#5629# => X"9ca00001",
		16#562a# => X"9ca00000",
		16#562b# => X"a4a500ff",
		16#562c# => X"bc250000",
		16#562d# => X"10000046",
		16#562e# => X"15000000",
		16#562f# => X"1840fff0",
		16#5630# => X"e0e31000",
		16#5631# => X"18407fdf",
		16#5632# => X"a842ffff",
		16#5633# => X"e4a71000",
		16#5634# => X"0c000039",
		16#5635# => X"9cc00001",
		16#5636# => X"a4c600ff",
		16#5637# => X"bc260000",
		16#5638# => X"1000003b",
		16#5639# => X"15000000",
		16#563a# => X"18408000",
		16#563b# => X"e0e31000",
		16#563c# => X"1840000f",
		16#563d# => X"a842ffff",
		16#563e# => X"e4a71000",
		16#563f# => X"0c000027",
		16#5640# => X"9ca00001",
		16#5641# => X"a4a500ff",
		16#5642# => X"bc250000",
		16#5643# => X"1000002c",
		16#5644# => X"15000000",
		16#5645# => X"1840000f",
		16#5646# => X"a842ffff",
		16#5647# => X"e4a31000",
		16#5648# => X"10000003",
		16#5649# => X"9cc00001",
		16#564a# => X"a8c50000",
		16#564b# => X"a4c600ff",
		16#564c# => X"bc260000",
		16#564d# => X"10000022",
		16#564e# => X"15000000",
		16#564f# => X"1840fff0",
		16#5650# => X"e0a31005",
		16#5651# => X"18407ff0",
		16#5652# => X"e1602802",
		16#5653# => X"e0631005",
		16#5654# => X"e0ab2804",
		16#5655# => X"e0c01802",
		16#5656# => X"e0661804",
		16#5657# => X"e1632803",
		16#5658# => X"ad6bffff",
		16#5659# => X"b96b005f",
		16#565a# => X"e1645803",
		16#565b# => X"9c210004",
		16#565c# => X"44004800",
		16#565d# => X"8441fffc",
		16#565e# => X"e0a31000",
		16#565f# => X"e0c02802",
		16#5660# => X"e0a62804",
		16#5661# => X"bd650000",
		16#5662# => X"0fffffc1",
		16#5663# => X"15000000",
		16#5664# => X"03fffff8",
		16#5665# => X"9c210004",
		16#5666# => X"a8a60000",
		16#5667# => X"a4a500ff",
		16#5668# => X"bc250000",
		16#5669# => X"0fffffdc",
		16#566a# => X"15000000",
		16#566b# => X"00000005",
		16#566c# => X"9c210004",
		16#566d# => X"03ffffc9",
		16#566e# => X"a8c50000",
		16#566f# => X"9c210004",
		16#5670# => X"9d600003",
		16#5671# => X"44004800",
		16#5672# => X"8441fffc",
		16#5673# => X"9c210004",
		16#5674# => X"9d600004",
		16#5675# => X"44004800",
		16#5676# => X"8441fffc",
		16#5677# => X"d7e117f8",
		16#5678# => X"a8440000",
		16#5679# => X"9884000e",
		16#567a# => X"d7e14ffc",
		16#567b# => X"0400068f",
		16#567c# => X"9c21fff8",
		16#567d# => X"bd8b0000",
		16#567e# => X"10000009",
		16#567f# => X"9c80efff",
		16#5680# => X"84620050",
		16#5681# => X"e0635800",
		16#5682# => X"d4021850",
		16#5683# => X"9c210008",
		16#5684# => X"8521fffc",
		16#5685# => X"44004800",
		16#5686# => X"8441fff8",
		16#5687# => X"9462000c",
		16#5688# => X"e0632003",
		16#5689# => X"dc02180c",
		16#568a# => X"9c210008",
		16#568b# => X"8521fffc",
		16#568c# => X"44004800",
		16#568d# => X"8441fff8",
		16#568e# => X"44004800",
		16#568f# => X"9d600000",
		16#5690# => X"d7e117ec",
		16#5691# => X"a8440000",
		16#5692# => X"9884000c",
		16#5693# => X"d7e177f0",
		16#5694# => X"d7e187f4",
		16#5695# => X"d7e197f8",
		16#5696# => X"d7e14ffc",
		16#5697# => X"a4e40100",
		16#5698# => X"9c21ffec",
		16#5699# => X"aa430000",
		16#569a# => X"aa050000",
		16#569b# => X"bc070000",
		16#569c# => X"10000007",
		16#569d# => X"a9c60000",
		16#569e# => X"9882000e",
		16#569f# => X"9ca00000",
		16#56a0# => X"0400064b",
		16#56a1# => X"9cc00002",
		16#56a2# => X"9882000c",
		16#56a3# => X"9ca0efff",
		16#56a4# => X"a8ce0000",
		16#56a5# => X"e0642803",
		16#56a6# => X"9882000e",
		16#56a7# => X"dc02180c",
		16#56a8# => X"9c210014",
		16#56a9# => X"a8720000",
		16#56aa# => X"a8b00000",
		16#56ab# => X"8521fffc",
		16#56ac# => X"8441ffec",
		16#56ad# => X"85c1fff0",
		16#56ae# => X"8601fff4",
		16#56af# => X"000004a9",
		16#56b0# => X"8641fff8",
		16#56b1# => X"d7e117f8",
		16#56b2# => X"a8440000",
		16#56b3# => X"9884000e",
		16#56b4# => X"d7e14ffc",
		16#56b5# => X"04000636",
		16#56b6# => X"9c21fff8",
		16#56b7# => X"bc2bffff",
		16#56b8# => X"0c00000a",
		16#56b9# => X"9c80efff",
		16#56ba# => X"9462000c",
		16#56bb# => X"a8631000",
		16#56bc# => X"d4025850",
		16#56bd# => X"dc02180c",
		16#56be# => X"9c210008",
		16#56bf# => X"8521fffc",
		16#56c0# => X"44004800",
		16#56c1# => X"8441fff8",
		16#56c2# => X"9462000c",
		16#56c3# => X"e0632003",
		16#56c4# => X"dc02180c",
		16#56c5# => X"9c210008",
		16#56c6# => X"8521fffc",
		16#56c7# => X"44004800",
		16#56c8# => X"8441fff8",
		16#56c9# => X"d7e14ffc",
		16#56ca# => X"9c21fffc",
		16#56cb# => X"9884000e",
		16#56cc# => X"9c210004",
		16#56cd# => X"8521fffc",
		16#56ce# => X"000004da",
		16#56cf# => X"15000000",
		16#56d0# => X"e1641804",
		16#56d1# => X"d7e117fc",
		16#56d2# => X"a56b0003",
		16#56d3# => X"bc2b0000",
		16#56d4# => X"10000024",
		16#56d5# => X"9c21fffc",
		16#56d6# => X"84a30000",
		16#56d7# => X"84c40000",
		16#56d8# => X"e4253000",
		16#56d9# => X"1000001f",
		16#56da# => X"1840fefe",
		16#56db# => X"a842feff",
		16#56dc# => X"e0c51000",
		16#56dd# => X"aca5ffff",
		16#56de# => X"18408080",
		16#56df# => X"e0a62803",
		16#56e0# => X"a8428080",
		16#56e1# => X"e0a51003",
		16#56e2# => X"bc250000",
		16#56e3# => X"0c00000b",
		16#56e4# => X"9c630004",
		16#56e5# => X"9c63fffc",
		16#56e6# => X"0000002a",
		16#56e7# => X"9c210004",
		16#56e8# => X"18408080",
		16#56e9# => X"a8428080",
		16#56ea# => X"e0c61003",
		16#56eb# => X"bc260000",
		16#56ec# => X"10000026",
		16#56ed# => X"9c630004",
		16#56ee# => X"1840fefe",
		16#56ef# => X"84a30000",
		16#56f0# => X"9c840004",
		16#56f1# => X"a842feff",
		16#56f2# => X"85040000",
		16#56f3# => X"e0e51000",
		16#56f4# => X"acc5ffff",
		16#56f5# => X"e4054000",
		16#56f6# => X"13fffff2",
		16#56f7# => X"e0c73003",
		16#56f8# => X"90a30000",
		16#56f9# => X"bc050000",
		16#56fa# => X"10000012",
		16#56fb# => X"15000000",
		16#56fc# => X"90c40000",
		16#56fd# => X"e4262800",
		16#56fe# => X"0c00000a",
		16#56ff# => X"9c630001",
		16#5700# => X"9c63ffff",
		16#5701# => X"0000000c",
		16#5702# => X"8d630000",
		16#5703# => X"90c40000",
		16#5704# => X"e4062800",
		16#5705# => X"0c000007",
		16#5706# => X"15000000",
		16#5707# => X"9c630001",
		16#5708# => X"90a30000",
		16#5709# => X"bc050000",
		16#570a# => X"0ffffff9",
		16#570b# => X"9c840001",
		16#570c# => X"8d630000",
		16#570d# => X"8c640000",
		16#570e# => X"e16b1802",
		16#570f# => X"9c210004",
		16#5710# => X"44004800",
		16#5711# => X"8441fffc",
		16#5712# => X"9c210004",
		16#5713# => X"9d600000",
		16#5714# => X"44004800",
		16#5715# => X"8441fffc",
		16#5716# => X"d7e197ec",
		16#5717# => X"d7e1a7f0",
		16#5718# => X"d7e1b7f4",
		16#5719# => X"d7e14ffc",
		16#571a# => X"d7e117e0",
		16#571b# => X"d7e177e4",
		16#571c# => X"d7e187e8",
		16#571d# => X"d7e1c7f8",
		16#571e# => X"85650008",
		16#571f# => X"9c21ffe0",
		16#5720# => X"aac50000",
		16#5721# => X"aa830000",
		16#5722# => X"bc2b0000",
		16#5723# => X"0c00002f",
		16#5724# => X"aa440000",
		16#5725# => X"84440064",
		16#5726# => X"a4422000",
		16#5727# => X"bc020000",
		16#5728# => X"1000002c",
		16#5729# => X"15000000",
		16#572a# => X"87050000",
		16#572b# => X"86180004",
		16#572c# => X"ba100042",
		16#572d# => X"bdb00000",
		16#572e# => X"1000001d",
		16#572f# => X"84580000",
		16#5730# => X"00000005",
		16#5731# => X"9dc00000",
		16#5732# => X"e5507000",
		16#5733# => X"0c000017",
		16#5734# => X"15000000",
		16#5735# => X"84820000",
		16#5736# => X"a8740000",
		16#5737# => X"a8b20000",
		16#5738# => X"040004eb",
		16#5739# => X"9dce0001",
		16#573a# => X"bc0bffff",
		16#573b# => X"0ffffff7",
		16#573c# => X"9c420004",
		16#573d# => X"9c400000",
		16#573e# => X"d4161008",
		16#573f# => X"d4161004",
		16#5740# => X"9c210020",
		16#5741# => X"8521fffc",
		16#5742# => X"8441ffe0",
		16#5743# => X"85c1ffe4",
		16#5744# => X"8601ffe8",
		16#5745# => X"8641ffec",
		16#5746# => X"8681fff0",
		16#5747# => X"86c1fff4",
		16#5748# => X"44004800",
		16#5749# => X"8701fff8",
		16#574a# => X"85760008",
		16#574b# => X"ba100002",
		16#574c# => X"e16b8002",
		16#574d# => X"bc0b0000",
		16#574e# => X"13ffffef",
		16#574f# => X"d4165808",
		16#5750# => X"03ffffdb",
		16#5751# => X"9f180008",
		16#5752# => X"03ffffee",
		16#5753# => X"d4055804",
		16#5754# => X"07fff427",
		16#5755# => X"9c400000",
		16#5756# => X"03ffffe9",
		16#5757# => X"d4161008",
		16#5758# => X"d7e177d8",
		16#5759# => X"d7e14ffc",
		16#575a# => X"d7e117d4",
		16#575b# => X"d7e187dc",
		16#575c# => X"d7e197e0",
		16#575d# => X"d7e1a7e4",
		16#575e# => X"d7e1b7e8",
		16#575f# => X"d7e1c7ec",
		16#5760# => X"d7e1d7f0",
		16#5761# => X"d7e1e7f4",
		16#5762# => X"d7e1f7f8",
		16#5763# => X"9c21fac4",
		16#5764# => X"a9c50000",
		16#5765# => X"d4011824",
		16#5766# => X"d4012020",
		16#5767# => X"bc030000",
		16#5768# => X"10000006",
		16#5769# => X"d4013014",
		16#576a# => X"84430038",
		16#576b# => X"bc220000",
		16#576c# => X"0c000335",
		16#576d# => X"15000000",
		16#576e# => X"84610020",
		16#576f# => X"9843000c",
		16#5770# => X"a4e2ffff",
		16#5771# => X"a4a72000",
		16#5772# => X"bc250000",
		16#5773# => X"1000000b",
		16#5774# => X"a4a70008",
		16#5775# => X"84a30064",
		16#5776# => X"9c60dfff",
		16#5777# => X"a8422000",
		16#5778# => X"84810020",
		16#5779# => X"e0a51803",
		16#577a# => X"dc04100c",
		16#577b# => X"d4042864",
		16#577c# => X"a4e2ffff",
		16#577d# => X"a4a70008",
		16#577e# => X"bc050000",
		16#577f# => X"100003b1",
		16#5780# => X"84810020",
		16#5781# => X"84a40010",
		16#5782# => X"bc250000",
		16#5783# => X"0c0003ae",
		16#5784# => X"84610024",
		16#5785# => X"a4e7001a",
		16#5786# => X"bc27000a",
		16#5787# => X"0c0002ed",
		16#5788# => X"84610020",
		16#5789# => X"9c400000",
		16#578a# => X"9c610500",
		16#578b# => X"9c8104ff",
		16#578c# => X"d4011804",
		16#578d# => X"d4011028",
		16#578e# => X"9c600000",
		16#578f# => X"9c410498",
		16#5790# => X"d4012000",
		16#5791# => X"d4011500",
		16#5792# => X"d4011d08",
		16#5793# => X"d4011d04",
		16#5794# => X"d401180c",
		16#5795# => X"aa420000",
		16#5796# => X"84610000",
		16#5797# => X"84410004",
		16#5798# => X"aace0000",
		16#5799# => X"e0421802",
		16#579a# => X"87410024",
		16#579b# => X"d401102c",
		16#579c# => X"87810020",
		16#579d# => X"90560000",
		16#579e# => X"aca20025",
		16#579f# => X"a4a500ff",
		16#57a0# => X"bc050000",
		16#57a1# => X"10000238",
		16#57a2# => X"15000000",
		16#57a3# => X"a44200ff",
		16#57a4# => X"bc020000",
		16#57a5# => X"10000234",
		16#57a6# => X"15000000",
		16#57a7# => X"00000005",
		16#57a8# => X"a8560000",
		16#57a9# => X"bc230000",
		16#57aa# => X"0c00000a",
		16#57ab# => X"e1c2b002",
		16#57ac# => X"9c420001",
		16#57ad# => X"90a20000",
		16#57ae# => X"ac650025",
		16#57af# => X"a46300ff",
		16#57b0# => X"bc030000",
		16#57b1# => X"0ffffff8",
		16#57b2# => X"a46500ff",
		16#57b3# => X"e1c2b002",
		16#57b4# => X"bc0e0000",
		16#57b5# => X"10000012",
		16#57b6# => X"bc050000",
		16#57b7# => X"84a10508",
		16#57b8# => X"84c10504",
		16#57b9# => X"e0a57000",
		16#57ba# => X"9cc60001",
		16#57bb# => X"d412b000",
		16#57bc# => X"d4127004",
		16#57bd# => X"d4012d08",
		16#57be# => X"bd460007",
		16#57bf# => X"1000028b",
		16#57c0# => X"d4013504",
		16#57c1# => X"9e520008",
		16#57c2# => X"8481000c",
		16#57c3# => X"e0847000",
		16#57c4# => X"d401200c",
		16#57c5# => X"90a20000",
		16#57c6# => X"bc050000",
		16#57c7# => X"1000021f",
		16#57c8# => X"9ca00000",
		16#57c9# => X"9ec20001",
		16#57ca# => X"9c400000",
		16#57cb# => X"9dc0ffff",
		16#57cc# => X"d801150f",
		16#57cd# => X"d4012810",
		16#57ce# => X"ab050000",
		16#57cf# => X"90d60000",
		16#57d0# => X"9ed60001",
		16#57d1# => X"9c46ffe0",
		16#57d2# => X"bc420058",
		16#57d3# => X"0c00004d",
		16#57d4# => X"18600001",
		16#57d5# => X"bc060000",
		16#57d6# => X"10000210",
		16#57d7# => X"d8012d0f",
		16#57d8# => X"9c600001",
		16#57d9# => X"9c800000",
		16#57da# => X"d4011808",
		16#57db# => X"d80134d8",
		16#57dc# => X"d801250f",
		16#57dd# => X"abc30000",
		16#57de# => X"9e0104d8",
		16#57df# => X"9c400000",
		16#57e0# => X"d4011018",
		16#57e1# => X"a4580002",
		16#57e2# => X"bc020000",
		16#57e3# => X"10000005",
		16#57e4# => X"a4980084",
		16#57e5# => X"84610008",
		16#57e6# => X"9c630002",
		16#57e7# => X"d4011808",
		16#57e8# => X"bc040000",
		16#57e9# => X"0c00014c",
		16#57ea# => X"d401201c",
		16#57eb# => X"84610010",
		16#57ec# => X"84810008",
		16#57ed# => X"e2832002",
		16#57ee# => X"bd540000",
		16#57ef# => X"0c000146",
		16#57f0# => X"bd540010",
		16#57f1# => X"0c000332",
		16#57f2# => X"15000000",
		16#57f3# => X"19c00001",
		16#57f4# => X"84a10508",
		16#57f5# => X"84c10504",
		16#57f6# => X"00000007",
		16#57f7# => X"a9ce8d9c",
		16#57f8# => X"9e520008",
		16#57f9# => X"9e94fff0",
		16#57fa# => X"bd540010",
		16#57fb# => X"0c00001a",
		16#57fc# => X"9d920008",
		16#57fd# => X"18600001",
		16#57fe# => X"9cc60001",
		16#57ff# => X"9ca50010",
		16#5800# => X"a8638d9c",
		16#5801# => X"9c800010",
		16#5802# => X"d4121800",
		16#5803# => X"d4122004",
		16#5804# => X"d4012d08",
		16#5805# => X"bd460007",
		16#5806# => X"0ffffff2",
		16#5807# => X"d4013504",
		16#5808# => X"a87a0000",
		16#5809# => X"a89c0000",
		16#580a# => X"07ffff0c",
		16#580b# => X"9ca10500",
		16#580c# => X"bc2b0000",
		16#580d# => X"100001e1",
		16#580e# => X"9e94fff0",
		16#580f# => X"9d8104a0",
		16#5810# => X"9e410498",
		16#5811# => X"84a10508",
		16#5812# => X"bd540010",
		16#5813# => X"13ffffea",
		16#5814# => X"84c10504",
		16#5815# => X"9cc60001",
		16#5816# => X"e0a5a000",
		16#5817# => X"d4127000",
		16#5818# => X"d412a004",
		16#5819# => X"d4012d08",
		16#581a# => X"bd460007",
		16#581b# => X"100002b9",
		16#581c# => X"d4013504",
		16#581d# => X"9dac0008",
		16#581e# => X"0000011a",
		16#581f# => X"aa4c0000",
		16#5820# => X"b8420002",
		16#5821# => X"a8638c28",
		16#5822# => X"e0421800",
		16#5823# => X"84420000",
		16#5824# => X"44001000",
		16#5825# => X"15000000",
		16#5826# => X"03ffffa9",
		16#5827# => X"ab180010",
		16#5828# => X"ab180010",
		16#5829# => X"a4b80010",
		16#582a# => X"bc050000",
		16#582b# => X"1000029e",
		16#582c# => X"a5180040",
		16#582d# => X"84610014",
		16#582e# => X"9ca00000",
		16#582f# => X"84430000",
		16#5830# => X"e1001002",
		16#5831# => X"9c630004",
		16#5832# => X"e1081004",
		16#5833# => X"d4011814",
		16#5834# => X"b908005f",
		16#5835# => X"9c600000",
		16#5836# => X"d8011d0f",
		16#5837# => X"bd8e0000",
		16#5838# => X"10000003",
		16#5839# => X"9c80ff7f",
		16#583a# => X"e3182003",
		16#583b# => X"e0c07002",
		16#583c# => X"e0c67004",
		16#583d# => X"bd860000",
		16#583e# => X"10000006",
		16#583f# => X"bc050001",
		16#5840# => X"bc080000",
		16#5841# => X"1000019b",
		16#5842# => X"bc250000",
		16#5843# => X"bc050001",
		16#5844# => X"10000270",
		16#5845# => X"bc050002",
		16#5846# => X"10000262",
		16#5847# => X"9e010500",
		16#5848# => X"a4a20007",
		16#5849# => X"9e10ffff",
		16#584a# => X"9ca50030",
		16#584b# => X"b8420043",
		16#584c# => X"bc220000",
		16#584d# => X"13fffffb",
		16#584e# => X"d8102800",
		16#584f# => X"a4580001",
		16#5850# => X"bc220000",
		16#5851# => X"0c000008",
		16#5852# => X"84410004",
		16#5853# => X"bc250030",
		16#5854# => X"0c0002d5",
		16#5855# => X"9c800030",
		16#5856# => X"9e10ffff",
		16#5857# => X"d8102000",
		16#5858# => X"84410004",
		16#5859# => X"e3c28002",
		16#585a# => X"d4017018",
		16#585b# => X"84810018",
		16#585c# => X"e57e2000",
		16#585d# => X"10000003",
		16#585e# => X"d401f008",
		16#585f# => X"d4012008",
		16#5860# => X"90c1050f",
		16#5861# => X"bc060000",
		16#5862# => X"13ffff7f",
		16#5863# => X"84410008",
		16#5864# => X"9c420001",
		16#5865# => X"03ffff7c",
		16#5866# => X"d4011008",
		16#5867# => X"ab180010",
		16#5868# => X"a4580010",
		16#5869# => X"bc020000",
		16#586a# => X"0c000009",
		16#586b# => X"84610014",
		16#586c# => X"a4580040",
		16#586d# => X"bc020000",
		16#586e# => X"10000005",
		16#586f# => X"84810014",
		16#5870# => X"9ca00001",
		16#5871# => X"0000025d",
		16#5872# => X"84440000",
		16#5873# => X"9ca00001",
		16#5874# => X"03ffffbc",
		16#5875# => X"84430000",
		16#5876# => X"84410014",
		16#5877# => X"84610014",
		16#5878# => X"84420000",
		16#5879# => X"9c630004",
		16#587a# => X"d4011010",
		16#587b# => X"bd620000",
		16#587c# => X"13ffff53",
		16#587d# => X"d4011814",
		16#587e# => X"e0401002",
		16#587f# => X"d4011010",
		16#5880# => X"03ffff4f",
		16#5881# => X"ab180004",
		16#5882# => X"03ffff4d",
		16#5883# => X"9ca0002b",
		16#5884# => X"03ffff4b",
		16#5885# => X"ab180080",
		16#5886# => X"90d60000",
		16#5887# => X"bc06002a",
		16#5888# => X"100002ba",
		16#5889# => X"9ed60001",
		16#588a# => X"9c46ffd0",
		16#588b# => X"bca20009",
		16#588c# => X"0c00000b",
		16#588d# => X"9dc00000",
		16#588e# => X"b88e0003",
		16#588f# => X"e1ce7000",
		16#5890# => X"90d60000",
		16#5891# => X"e1ce2000",
		16#5892# => X"e1ce1000",
		16#5893# => X"9c46ffd0",
		16#5894# => X"bca20009",
		16#5895# => X"13fffff9",
		16#5896# => X"9ed60001",
		16#5897# => X"bd6e0000",
		16#5898# => X"13ffff3a",
		16#5899# => X"9c46ffe0",
		16#589a# => X"03ffff38",
		16#589b# => X"9dc0ffff",
		16#589c# => X"a4580010",
		16#589d# => X"bc020000",
		16#589e# => X"0c00024a",
		16#589f# => X"d8012d0f",
		16#58a0# => X"a4580040",
		16#58a1# => X"bc020000",
		16#58a2# => X"10000247",
		16#58a3# => X"84610014",
		16#58a4# => X"8481000c",
		16#58a5# => X"84430000",
		16#58a6# => X"9c630004",
		16#58a7# => X"d4011814",
		16#58a8# => X"03fffef5",
		16#58a9# => X"dc022000",
		16#58aa# => X"18800001",
		16#58ab# => X"d8012d0f",
		16#58ac# => X"a88488b7",
		16#58ad# => X"d4012028",
		16#58ae# => X"a4580010",
		16#58af# => X"bc020000",
		16#58b0# => X"0c000007",
		16#58b1# => X"84610014",
		16#58b2# => X"a4580040",
		16#58b3# => X"bc020000",
		16#58b4# => X"0c00023e",
		16#58b5# => X"84810014",
		16#58b6# => X"84610014",
		16#58b7# => X"84430000",
		16#58b8# => X"9c630004",
		16#58b9# => X"d4011814",
		16#58ba# => X"e1001002",
		16#58bb# => X"e1081004",
		16#58bc# => X"b908005f",
		16#58bd# => X"bc080000",
		16#58be# => X"13ffff77",
		16#58bf# => X"9ca00002",
		16#58c0# => X"a4b80001",
		16#58c1# => X"bc050000",
		16#58c2# => X"10000008",
		16#58c3# => X"9c800030",
		16#58c4# => X"d801350d",
		16#58c5# => X"d801250c",
		16#58c6# => X"ab180002",
		16#58c7# => X"9d000001",
		16#58c8# => X"03ffff6d",
		16#58c9# => X"9ca00002",
		16#58ca# => X"03ffff6b",
		16#58cb# => X"9ca00002",
		16#58cc# => X"84810014",
		16#58cd# => X"9c600030",
		16#58ce# => X"84440000",
		16#58cf# => X"9c800078",
		16#58d0# => X"e1001002",
		16#58d1# => X"d8011d0c",
		16#58d2# => X"d801250d",
		16#58d3# => X"84610014",
		16#58d4# => X"18800001",
		16#58d5# => X"e1081004",
		16#58d6# => X"9c630004",
		16#58d7# => X"a88488b7",
		16#58d8# => X"ab180002",
		16#58d9# => X"b908005f",
		16#58da# => X"d4011814",
		16#58db# => X"d4012028",
		16#58dc# => X"03ffff59",
		16#58dd# => X"9ca00002",
		16#58de# => X"84410014",
		16#58df# => X"9c600000",
		16#58e0# => X"9c820004",
		16#58e1# => X"d8011d0f",
		16#58e2# => X"d4012014",
		16#58e3# => X"86020000",
		16#58e4# => X"bc300000",
		16#58e5# => X"0c000233",
		16#58e6# => X"bd8e0000",
		16#58e7# => X"1000022c",
		16#58e8# => X"a8700000",
		16#58e9# => X"9c800000",
		16#58ea# => X"07fff521",
		16#58eb# => X"a8ae0000",
		16#58ec# => X"bc0b0000",
		16#58ed# => X"10000251",
		16#58ee# => X"abce0000",
		16#58ef# => X"e3cb8002",
		16#58f0# => X"e55e7000",
		16#58f1# => X"0c000220",
		16#58f2# => X"9c400000",
		16#58f3# => X"9c600000",
		16#58f4# => X"abce0000",
		16#58f5# => X"03ffff66",
		16#58f6# => X"d4011818",
		16#58f7# => X"03fffed8",
		16#58f8# => X"ab180001",
		16#58f9# => X"bc250000",
		16#58fa# => X"13fffed5",
		16#58fb# => X"15000000",
		16#58fc# => X"03fffed3",
		16#58fd# => X"9ca00020",
		16#58fe# => X"03fffed1",
		16#58ff# => X"ab180040",
		16#5900# => X"d8012d0f",
		16#5901# => X"a4580010",
		16#5902# => X"bc020000",
		16#5903# => X"0c000007",
		16#5904# => X"84610014",
		16#5905# => X"a4580040",
		16#5906# => X"bc020000",
		16#5907# => X"0c0001f0",
		16#5908# => X"84810014",
		16#5909# => X"84610014",
		16#590a# => X"84430000",
		16#590b# => X"9c630004",
		16#590c# => X"bd820000",
		16#590d# => X"100001ef",
		16#590e# => X"d4011814",
		16#590f# => X"e1001002",
		16#5910# => X"9ca00001",
		16#5911# => X"e1081004",
		16#5912# => X"03ffff25",
		16#5913# => X"b908005f",
		16#5914# => X"84410014",
		16#5915# => X"9c600001",
		16#5916# => X"84a20000",
		16#5917# => X"9c800000",
		16#5918# => X"9c420004",
		16#5919# => X"d4011808",
		16#591a# => X"d8012cd8",
		16#591b# => X"d801250f",
		16#591c# => X"d4011014",
		16#591d# => X"abc30000",
		16#591e# => X"03fffec1",
		16#591f# => X"9e0104d8",
		16#5920# => X"18800001",
		16#5921# => X"d8012d0f",
		16#5922# => X"a88488a6",
		16#5923# => X"03ffff8b",
		16#5924# => X"d4012028",
		16#5925# => X"d8012d0f",
		16#5926# => X"03ffffdb",
		16#5927# => X"ab180010",
		16#5928# => X"9c600000",
		16#5929# => X"9c46ffd0",
		16#592a# => X"b8830003",
		16#592b# => X"e0631800",
		16#592c# => X"90d60000",
		16#592d# => X"e0632000",
		16#592e# => X"e0621800",
		16#592f# => X"9c46ffd0",
		16#5930# => X"bca20009",
		16#5931# => X"13fffff9",
		16#5932# => X"9ed60001",
		16#5933# => X"03fffe9e",
		16#5934# => X"d4011810",
		16#5935# => X"9db20008",
		16#5936# => X"84a10508",
		16#5937# => X"84c10504",
		16#5938# => X"9181050f",
		16#5939# => X"bc0c0000",
		16#593a# => X"1000000f",
		16#593b# => X"bc020000",
		16#593c# => X"9cc60001",
		16#593d# => X"9ca50001",
		16#593e# => X"9c61050f",
		16#593f# => X"9c800001",
		16#5940# => X"d4121800",
		16#5941# => X"d4122004",
		16#5942# => X"d4012d08",
		16#5943# => X"bd460007",
		16#5944# => X"1000011a",
		16#5945# => X"d4013504",
		16#5946# => X"aa4d0000",
		16#5947# => X"9dad0008",
		16#5948# => X"bc020000",
		16#5949# => X"1000000f",
		16#594a# => X"8481001c",
		16#594b# => X"9cc60001",
		16#594c# => X"9ca50002",
		16#594d# => X"9c41050c",
		16#594e# => X"9c600002",
		16#594f# => X"d4121000",
		16#5950# => X"d4121804",
		16#5951# => X"d4012d08",
		16#5952# => X"bd460007",
		16#5953# => X"10000116",
		16#5954# => X"d4013504",
		16#5955# => X"aa4d0000",
		16#5956# => X"9dad0008",
		16#5957# => X"8481001c",
		16#5958# => X"bc240080",
		16#5959# => X"0c0000ab",
		16#595a# => X"84410010",
		16#595b# => X"84810018",
		16#595c# => X"e1c4f002",
		16#595d# => X"bdae0000",
		16#595e# => X"1000002e",
		16#595f# => X"bdae0010",
		16#5960# => X"100001ad",
		16#5961# => X"15000000",
		16#5962# => X"18400001",
		16#5963# => X"00000007",
		16#5964# => X"a8428d8c",
		16#5965# => X"9e520008",
		16#5966# => X"9dcefff0",
		16#5967# => X"bd4e0010",
		16#5968# => X"0c00001a",
		16#5969# => X"9d920008",
		16#596a# => X"18600001",
		16#596b# => X"9cc60001",
		16#596c# => X"9ca50010",
		16#596d# => X"a8638d8c",
		16#596e# => X"9c800010",
		16#596f# => X"d4121800",
		16#5970# => X"d4122004",
		16#5971# => X"d4012d08",
		16#5972# => X"bd460007",
		16#5973# => X"0ffffff2",
		16#5974# => X"d4013504",
		16#5975# => X"a87a0000",
		16#5976# => X"a89c0000",
		16#5977# => X"07fffd9f",
		16#5978# => X"9ca10500",
		16#5979# => X"bc2b0000",
		16#597a# => X"10000074",
		16#597b# => X"9dcefff0",
		16#597c# => X"9d8104a0",
		16#597d# => X"9e410498",
		16#597e# => X"84a10508",
		16#597f# => X"bd4e0010",
		16#5980# => X"13ffffea",
		16#5981# => X"84c10504",
		16#5982# => X"9cc60001",
		16#5983# => X"e0a57000",
		16#5984# => X"d4121000",
		16#5985# => X"d4127004",
		16#5986# => X"d4012d08",
		16#5987# => X"bd460007",
		16#5988# => X"100000cb",
		16#5989# => X"d4013504",
		16#598a# => X"9dac0008",
		16#598b# => X"aa4c0000",
		16#598c# => X"9cc60001",
		16#598d# => X"e0a5f000",
		16#598e# => X"d4128000",
		16#598f# => X"d412f004",
		16#5990# => X"d4012d08",
		16#5991# => X"bda60007",
		16#5992# => X"0c0000a4",
		16#5993# => X"d4013504",
		16#5994# => X"a4d80004",
		16#5995# => X"bc260000",
		16#5996# => X"0c000032",
		16#5997# => X"84410008",
		16#5998# => X"84610010",
		16#5999# => X"84810008",
		16#599a# => X"e0432002",
		16#599b# => X"bd420000",
		16#599c# => X"0c00002b",
		16#599d# => X"bda20010",
		16#599e# => X"1000018e",
		16#599f# => X"15000000",
		16#59a0# => X"19c00001",
		16#59a1# => X"84c10504",
		16#59a2# => X"00000006",
		16#59a3# => X"a9ce8d9c",
		16#59a4# => X"9c42fff0",
		16#59a5# => X"bd420010",
		16#59a6# => X"0c000019",
		16#59a7# => X"9dad0008",
		16#59a8# => X"18600001",
		16#59a9# => X"9cc60001",
		16#59aa# => X"9ca50010",
		16#59ab# => X"a8638d9c",
		16#59ac# => X"9c800010",
		16#59ad# => X"d40d1800",
		16#59ae# => X"d40d2004",
		16#59af# => X"d4012d08",
		16#59b0# => X"bd460007",
		16#59b1# => X"0ffffff3",
		16#59b2# => X"d4013504",
		16#59b3# => X"a87a0000",
		16#59b4# => X"a89c0000",
		16#59b5# => X"07fffd61",
		16#59b6# => X"9ca10500",
		16#59b7# => X"bc2b0000",
		16#59b8# => X"10000036",
		16#59b9# => X"9c42fff0",
		16#59ba# => X"9da10498",
		16#59bb# => X"84a10508",
		16#59bc# => X"bd420010",
		16#59bd# => X"13ffffeb",
		16#59be# => X"84c10504",
		16#59bf# => X"9cc60001",
		16#59c0# => X"e0a22800",
		16#59c1# => X"d40d7000",
		16#59c2# => X"d40d1004",
		16#59c3# => X"d4012d08",
		16#59c4# => X"bda60007",
		16#59c5# => X"0c00011a",
		16#59c6# => X"d4013504",
		16#59c7# => X"84410008",
		16#59c8# => X"84610010",
		16#59c9# => X"e5621800",
		16#59ca# => X"10000003",
		16#59cb# => X"8481000c",
		16#59cc# => X"a8430000",
		16#59cd# => X"bc050000",
		16#59ce# => X"e0841000",
		16#59cf# => X"0c000070",
		16#59d0# => X"d401200c",
		16#59d1# => X"9c400000",
		16#59d2# => X"d4011504",
		16#59d3# => X"90560000",
		16#59d4# => X"aca20025",
		16#59d5# => X"a4a500ff",
		16#59d6# => X"bc050000",
		16#59d7# => X"0ffffdcc",
		16#59d8# => X"9e410498",
		16#59d9# => X"a8560000",
		16#59da# => X"03fffdec",
		16#59db# => X"90b60000",
		16#59dc# => X"1000006c",
		16#59dd# => X"abc80000",
		16#59de# => X"a4580001",
		16#59df# => X"bc020000",
		16#59e0# => X"100000c5",
		16#59e1# => X"9c400030",
		16#59e2# => X"87c1002c",
		16#59e3# => X"d80114ff",
		16#59e4# => X"03fffe76",
		16#59e5# => X"9e0104ff",
		16#59e6# => X"84410508",
		16#59e7# => X"bc020000",
		16#59e8# => X"10000007",
		16#59e9# => X"84610020",
		16#59ea# => X"84610024",
		16#59eb# => X"84810020",
		16#59ec# => X"07fffd2a",
		16#59ed# => X"9ca10500",
		16#59ee# => X"84610020",
		16#59ef# => X"9443000c",
		16#59f0# => X"a4420040",
		16#59f1# => X"bc020000",
		16#59f2# => X"10000005",
		16#59f3# => X"8561000c",
		16#59f4# => X"9c80ffff",
		16#59f5# => X"d401200c",
		16#59f6# => X"8561000c",
		16#59f7# => X"9c21053c",
		16#59f8# => X"8521fffc",
		16#59f9# => X"8441ffd4",
		16#59fa# => X"85c1ffd8",
		16#59fb# => X"8601ffdc",
		16#59fc# => X"8641ffe0",
		16#59fd# => X"8681ffe4",
		16#59fe# => X"86c1ffe8",
		16#59ff# => X"8701ffec",
		16#5a00# => X"8741fff0",
		16#5a01# => X"8781fff4",
		16#5a02# => X"44004800",
		16#5a03# => X"87c1fff8",
		16#5a04# => X"84610008",
		16#5a05# => X"e2821802",
		16#5a06# => X"bd540000",
		16#5a07# => X"0c0000f9",
		16#5a08# => X"bdb40010",
		16#5a09# => X"10000131",
		16#5a0a# => X"15000000",
		16#5a0b# => X"18400001",
		16#5a0c# => X"00000007",
		16#5a0d# => X"a8428d8c",
		16#5a0e# => X"9e520008",
		16#5a0f# => X"9e94fff0",
		16#5a10# => X"bd540010",
		16#5a11# => X"0c00001a",
		16#5a12# => X"9d920008",
		16#5a13# => X"18800001",
		16#5a14# => X"9cc60001",
		16#5a15# => X"9ca50010",
		16#5a16# => X"a8848d8c",
		16#5a17# => X"9c600010",
		16#5a18# => X"d4122000",
		16#5a19# => X"d4121804",
		16#5a1a# => X"d4012d08",
		16#5a1b# => X"bd460007",
		16#5a1c# => X"0ffffff2",
		16#5a1d# => X"d4013504",
		16#5a1e# => X"a87a0000",
		16#5a1f# => X"a89c0000",
		16#5a20# => X"07fffcf6",
		16#5a21# => X"9ca10500",
		16#5a22# => X"bc2b0000",
		16#5a23# => X"13ffffcb",
		16#5a24# => X"9e94fff0",
		16#5a25# => X"9d8104a0",
		16#5a26# => X"9e410498",
		16#5a27# => X"84a10508",
		16#5a28# => X"bd540010",
		16#5a29# => X"13ffffea",
		16#5a2a# => X"84c10504",
		16#5a2b# => X"9cc60001",
		16#5a2c# => X"e0a5a000",
		16#5a2d# => X"d4121000",
		16#5a2e# => X"d412a004",
		16#5a2f# => X"d4012d08",
		16#5a30# => X"bd460007",
		16#5a31# => X"100000d1",
		16#5a32# => X"d4013504",
		16#5a33# => X"9dac0008",
		16#5a34# => X"03ffff27",
		16#5a35# => X"aa4c0000",
		16#5a36# => X"a87a0000",
		16#5a37# => X"a89c0000",
		16#5a38# => X"07fffcde",
		16#5a39# => X"9ca10500",
		16#5a3a# => X"bc2b0000",
		16#5a3b# => X"13ffffb3",
		16#5a3c# => X"9da10498",
		16#5a3d# => X"03ffff57",
		16#5a3e# => X"84a10508",
		16#5a3f# => X"a87a0000",
		16#5a40# => X"a89c0000",
		16#5a41# => X"07fffcd5",
		16#5a42# => X"9ca10500",
		16#5a43# => X"bc2b0000",
		16#5a44# => X"0fffff8e",
		16#5a45# => X"9c400000",
		16#5a46# => X"03ffffa9",
		16#5a47# => X"84610020",
		16#5a48# => X"03fffe12",
		16#5a49# => X"9e010500",
		16#5a4a# => X"a87a0000",
		16#5a4b# => X"a89c0000",
		16#5a4c# => X"07fffcca",
		16#5a4d# => X"9ca10500",
		16#5a4e# => X"bc2b0000",
		16#5a4f# => X"13ffff9f",
		16#5a50# => X"9e410498",
		16#5a51# => X"03fffd72",
		16#5a52# => X"8481000c",
		16#5a53# => X"a87a0000",
		16#5a54# => X"a89c0000",
		16#5a55# => X"07fffcc1",
		16#5a56# => X"9ca10500",
		16#5a57# => X"bc2b0000",
		16#5a58# => X"13ffff96",
		16#5a59# => X"9da104a0",
		16#5a5a# => X"9e410498",
		16#5a5b# => X"84a10508",
		16#5a5c# => X"03ffff30",
		16#5a5d# => X"84c10504",
		16#5a5e# => X"a87a0000",
		16#5a5f# => X"a89c0000",
		16#5a60# => X"07fffcb6",
		16#5a61# => X"9ca10500",
		16#5a62# => X"bc2b0000",
		16#5a63# => X"13ffff8b",
		16#5a64# => X"9da104a0",
		16#5a65# => X"9e410498",
		16#5a66# => X"84a10508",
		16#5a67# => X"03fffee1",
		16#5a68# => X"84c10504",
		16#5a69# => X"a87a0000",
		16#5a6a# => X"a89c0000",
		16#5a6b# => X"07fffcab",
		16#5a6c# => X"9ca10500",
		16#5a6d# => X"bc2b0000",
		16#5a6e# => X"13ffff80",
		16#5a6f# => X"9da104a0",
		16#5a70# => X"9e410498",
		16#5a71# => X"84a10508",
		16#5a72# => X"03fffee5",
		16#5a73# => X"84c10504",
		16#5a74# => X"98e3000e",
		16#5a75# => X"bd870000",
		16#5a76# => X"13fffd13",
		16#5a77# => X"9c80fffd",
		16#5a78# => X"9e010430",
		16#5a79# => X"e0422003",
		16#5a7a# => X"85e30064",
		16#5a7b# => X"85a3001c",
		16#5a7c# => X"85830024",
		16#5a7d# => X"9d610030",
		16#5a7e# => X"9d000400",
		16#5a7f# => X"dc01143c",
		16#5a80# => X"84610024",
		16#5a81# => X"9c400000",
		16#5a82# => X"a8900000",
		16#5a83# => X"a8ae0000",
		16#5a84# => X"84c10014",
		16#5a85# => X"d4017c94",
		16#5a86# => X"dc013c3e",
		16#5a87# => X"d4016c4c",
		16#5a88# => X"d4016454",
		16#5a89# => X"d4015c30",
		16#5a8a# => X"d4015c40",
		16#5a8b# => X"d4014438",
		16#5a8c# => X"d4014444",
		16#5a8d# => X"07fffccb",
		16#5a8e# => X"d4011448",
		16#5a8f# => X"e58b1000",
		16#5a90# => X"10000008",
		16#5a91# => X"d401580c",
		16#5a92# => X"84610024",
		16#5a93# => X"07ffeded",
		16#5a94# => X"a8900000",
		16#5a95# => X"e42b1000",
		16#5a96# => X"100000aa",
		16#5a97# => X"9c60ffff",
		16#5a98# => X"9441043c",
		16#5a99# => X"a4420040",
		16#5a9a# => X"bc020000",
		16#5a9b# => X"13ffff5b",
		16#5a9c# => X"84810020",
		16#5a9d# => X"9444000c",
		16#5a9e# => X"a8420040",
		16#5a9f# => X"03ffff57",
		16#5aa0# => X"dc04100c",
		16#5aa1# => X"07ffeeed",
		16#5aa2# => X"15000000",
		16#5aa3# => X"03fffccc",
		16#5aa4# => X"84610020",
		16#5aa5# => X"abc50000",
		16#5aa6# => X"03fffdb4",
		16#5aa7# => X"9e010500",
		16#5aa8# => X"84810028",
		16#5aa9# => X"a462000f",
		16#5aaa# => X"9e10ffff",
		16#5aab# => X"e0641800",
		16#5aac# => X"b8420044",
		16#5aad# => X"8c630000",
		16#5aae# => X"bc220000",
		16#5aaf# => X"13fffffa",
		16#5ab0# => X"d8101800",
		16#5ab1# => X"84810004",
		16#5ab2# => X"03fffda8",
		16#5ab3# => X"e3c48002",
		16#5ab4# => X"bc420009",
		16#5ab5# => X"0c00000e",
		16#5ab6# => X"9e010500",
		16#5ab7# => X"a8620000",
		16#5ab8# => X"9c80000a",
		16#5ab9# => X"040004b7",
		16#5aba# => X"9e10ffff",
		16#5abb# => X"9d6b0030",
		16#5abc# => X"a8620000",
		16#5abd# => X"9c80000a",
		16#5abe# => X"07ffcb0e",
		16#5abf# => X"d8105800",
		16#5ac0# => X"bc4b0009",
		16#5ac1# => X"13fffff6",
		16#5ac2# => X"a84b0000",
		16#5ac3# => X"9e10ffff",
		16#5ac4# => X"84610004",
		16#5ac5# => X"9c420030",
		16#5ac6# => X"e3c38002",
		16#5ac7# => X"03fffd93",
		16#5ac8# => X"d8101000",
		16#5ac9# => X"bc080000",
		16#5aca# => X"10000025",
		16#5acb# => X"84610014",
		16#5acc# => X"84810014",
		16#5acd# => X"84440000",
		16#5ace# => X"a442ffff",
		16#5acf# => X"9c840004",
		16#5ad0# => X"e1001002",
		16#5ad1# => X"d4012014",
		16#5ad2# => X"03fffd63",
		16#5ad3# => X"b908005f",
		16#5ad4# => X"a87a0000",
		16#5ad5# => X"a89c0000",
		16#5ad6# => X"07fffc40",
		16#5ad7# => X"9ca10500",
		16#5ad8# => X"bc2b0000",
		16#5ad9# => X"13ffff15",
		16#5ada# => X"9da104a0",
		16#5adb# => X"9e410498",
		16#5adc# => X"84a10508",
		16#5add# => X"03fffe5b",
		16#5ade# => X"84c10504",
		16#5adf# => X"a87a0000",
		16#5ae0# => X"a89c0000",
		16#5ae1# => X"07fffc35",
		16#5ae2# => X"9ca10500",
		16#5ae3# => X"bc2b0000",
		16#5ae4# => X"13ffff0b",
		16#5ae5# => X"84610020",
		16#5ae6# => X"03fffee1",
		16#5ae7# => X"84a10508",
		16#5ae8# => X"84610014",
		16#5ae9# => X"8481000c",
		16#5aea# => X"84430000",
		16#5aeb# => X"9c630004",
		16#5aec# => X"d4011814",
		16#5aed# => X"03fffcb0",
		16#5aee# => X"d4022000",
		16#5aef# => X"a8a80000",
		16#5af0# => X"03fffd40",
		16#5af1# => X"84430000",
		16#5af2# => X"84440000",
		16#5af3# => X"9c840004",
		16#5af4# => X"a442ffff",
		16#5af5# => X"03fffdc5",
		16#5af6# => X"d4012014",
		16#5af7# => X"98440002",
		16#5af8# => X"9c840004",
		16#5af9# => X"bd820000",
		16#5afa# => X"0ffffe15",
		16#5afb# => X"d4012014",
		16#5afc# => X"9c80002d",
		16#5afd# => X"e0401002",
		16#5afe# => X"03fffe11",
		16#5aff# => X"d801250f",
		16#5b00# => X"03fffe5b",
		16#5b01# => X"9db20008",
		16#5b02# => X"a87a0000",
		16#5b03# => X"a89c0000",
		16#5b04# => X"07fffc12",
		16#5b05# => X"9ca10500",
		16#5b06# => X"bc2b0000",
		16#5b07# => X"13fffee7",
		16#5b08# => X"9da104a0",
		16#5b09# => X"9e410498",
		16#5b0a# => X"84a10508",
		16#5b0b# => X"03fffe50",
		16#5b0c# => X"84c10504",
		16#5b0d# => X"18400001",
		16#5b0e# => X"a98d0000",
		16#5b0f# => X"03fffe73",
		16#5b10# => X"a8428d8c",
		16#5b11# => X"03fffd4a",
		16#5b12# => X"d4011018",
		16#5b13# => X"9c400000",
		16#5b14# => X"07ffdb74",
		16#5b15# => X"d4011018",
		16#5b16# => X"03fffd45",
		16#5b17# => X"abcb0000",
		16#5b18# => X"bcae0006",
		16#5b19# => X"10000003",
		16#5b1a# => X"abce0000",
		16#5b1b# => X"9fc00006",
		16#5b1c# => X"ac5effff",
		16#5b1d# => X"1a000001",
		16#5b1e# => X"b842009f",
		16#5b1f# => X"aa1088c8",
		16#5b20# => X"e05e1003",
		16#5b21# => X"03fffcbe",
		16#5b22# => X"d4011008",
		16#5b23# => X"19c00001",
		16#5b24# => X"9d920008",
		16#5b25# => X"84a10508",
		16#5b26# => X"84c10504",
		16#5b27# => X"03fffcee",
		16#5b28# => X"a9ce8d9c",
		16#5b29# => X"84610004",
		16#5b2a# => X"03fffd30",
		16#5b2b# => X"e3c38002",
		16#5b2c# => X"19c00001",
		16#5b2d# => X"84c10504",
		16#5b2e# => X"03fffe91",
		16#5b2f# => X"a9ce8d9c",
		16#5b30# => X"84610024",
		16#5b31# => X"9c40ffff",
		16#5b32# => X"07ffe454",
		16#5b33# => X"d401100c",
		16#5b34# => X"bc2b0000",
		16#5b35# => X"13fffec1",
		16#5b36# => X"84610020",
		16#5b37# => X"9843000c",
		16#5b38# => X"03fffc4d",
		16#5b39# => X"a4e2ffff",
		16#5b3a# => X"18400001",
		16#5b3b# => X"a98d0000",
		16#5b3c# => X"03fffeef",
		16#5b3d# => X"a8428d8c",
		16#5b3e# => X"03fffd1d",
		16#5b3f# => X"d4015818",
		16#5b40# => X"03ffff58",
		16#5b41# => X"d401180c",
		16#5b42# => X"84810014",
		16#5b43# => X"85c40000",
		16#5b44# => X"bd8e0000",
		16#5b45# => X"10000004",
		16#5b46# => X"9c440004",
		16#5b47# => X"03fffc88",
		16#5b48# => X"d4011014",
		16#5b49# => X"d4011014",
		16#5b4a# => X"03fffc85",
		16#5b4b# => X"9dc0ffff",
		16#5b4c# => X"a8e40000",
		16#5b4d# => X"a8830000",
		16#5b4e# => X"18600001",
		16#5b4f# => X"d7e14ffc",
		16#5b50# => X"a863ade4",
		16#5b51# => X"9c21fffc",
		16#5b52# => X"84630000",
		16#5b53# => X"9c210004",
		16#5b54# => X"a8c50000",
		16#5b55# => X"8521fffc",
		16#5b56# => X"03fffc02",
		16#5b57# => X"a8a70000",
		16#5b58# => X"d7e117f4",
		16#5b59# => X"18400001",
		16#5b5a# => X"d7e177f8",
		16#5b5b# => X"a842c508",
		16#5b5c# => X"a9c30000",
		16#5b5d# => X"a8640000",
		16#5b5e# => X"a8850000",
		16#5b5f# => X"a8a60000",
		16#5b60# => X"9cc00000",
		16#5b61# => X"d7e14ffc",
		16#5b62# => X"d4023000",
		16#5b63# => X"040003cf",
		16#5b64# => X"9c21fff4",
		16#5b65# => X"bc2bffff",
		16#5b66# => X"0c000007",
		16#5b67# => X"15000000",
		16#5b68# => X"9c21000c",
		16#5b69# => X"8521fffc",
		16#5b6a# => X"8441fff4",
		16#5b6b# => X"44004800",
		16#5b6c# => X"85c1fff8",
		16#5b6d# => X"84420000",
		16#5b6e# => X"bc020000",
		16#5b6f# => X"13fffff9",
		16#5b70# => X"15000000",
		16#5b71# => X"d40e1000",
		16#5b72# => X"9c21000c",
		16#5b73# => X"8521fffc",
		16#5b74# => X"8441fff4",
		16#5b75# => X"44004800",
		16#5b76# => X"85c1fff8",
		16#5b77# => X"e0852306",
		16#5b78# => X"d7e117f8",
		16#5b79# => X"d7e14ffc",
		16#5b7a# => X"07ffd610",
		16#5b7b# => X"9c21fff8",
		16#5b7c# => X"bc0b0000",
		16#5b7d# => X"1000001e",
		16#5b7e# => X"a84b0000",
		16#5b7f# => X"9c60fffc",
		16#5b80# => X"84abfffc",
		16#5b81# => X"e0a51803",
		16#5b82# => X"e0a51800",
		16#5b83# => X"bc450024",
		16#5b84# => X"1000001c",
		16#5b85# => X"bca50013",
		16#5b86# => X"10000010",
		16#5b87# => X"a86b0000",
		16#5b88# => X"9c800000",
		16#5b89# => X"9c6b0008",
		16#5b8a# => X"d40b2000",
		16#5b8b# => X"bca5001b",
		16#5b8c# => X"1000000a",
		16#5b8d# => X"d40b2004",
		16#5b8e# => X"d4032000",
		16#5b8f# => X"d40b200c",
		16#5b90# => X"bc250024",
		16#5b91# => X"10000005",
		16#5b92# => X"9c6b0010",
		16#5b93# => X"d4032000",
		16#5b94# => X"d40b2014",
		16#5b95# => X"9c6b0018",
		16#5b96# => X"9ca00000",
		16#5b97# => X"9c830004",
		16#5b98# => X"d4032800",
		16#5b99# => X"d4042800",
		16#5b9a# => X"d4042804",
		16#5b9b# => X"9c210008",
		16#5b9c# => X"a9620000",
		16#5b9d# => X"8521fffc",
		16#5b9e# => X"44004800",
		16#5b9f# => X"8441fff8",
		16#5ba0# => X"a86b0000",
		16#5ba1# => X"07fff358",
		16#5ba2# => X"9c800000",
		16#5ba3# => X"9c210008",
		16#5ba4# => X"a9620000",
		16#5ba5# => X"8521fffc",
		16#5ba6# => X"44004800",
		16#5ba7# => X"8441fff8",
		16#5ba8# => X"d7e117f4",
		16#5ba9# => X"18400001",
		16#5baa# => X"d7e177f8",
		16#5bab# => X"a842c508",
		16#5bac# => X"a9c30000",
		16#5bad# => X"a8640000",
		16#5bae# => X"9c800000",
		16#5baf# => X"d7e14ffc",
		16#5bb0# => X"d4022000",
		16#5bb1# => X"0400020e",
		16#5bb2# => X"9c21fff4",
		16#5bb3# => X"bc2bffff",
		16#5bb4# => X"0c000007",
		16#5bb5# => X"15000000",
		16#5bb6# => X"9c21000c",
		16#5bb7# => X"8521fffc",
		16#5bb8# => X"8441fff4",
		16#5bb9# => X"44004800",
		16#5bba# => X"85c1fff8",
		16#5bbb# => X"84420000",
		16#5bbc# => X"bc020000",
		16#5bbd# => X"13fffff9",
		16#5bbe# => X"15000000",
		16#5bbf# => X"d40e1000",
		16#5bc0# => X"9c21000c",
		16#5bc1# => X"8521fffc",
		16#5bc2# => X"8441fff4",
		16#5bc3# => X"44004800",
		16#5bc4# => X"85c1fff8",
		16#5bc5# => X"d7e117f0",
		16#5bc6# => X"d7e177f4",
		16#5bc7# => X"d7e187f8",
		16#5bc8# => X"d7e14ffc",
		16#5bc9# => X"a8440000",
		16#5bca# => X"9c21fff0",
		16#5bcb# => X"a9c30000",
		16#5bcc# => X"bc040000",
		16#5bcd# => X"10000037",
		16#5bce# => X"aa040000",
		16#5bcf# => X"07ffee74",
		16#5bd0# => X"15000000",
		16#5bd1# => X"bc0e0000",
		16#5bd2# => X"10000006",
		16#5bd3# => X"15000000",
		16#5bd4# => X"846e0038",
		16#5bd5# => X"bc230000",
		16#5bd6# => X"0c000035",
		16#5bd7# => X"15000000",
		16#5bd8# => X"9a02000c",
		16#5bd9# => X"bc300000",
		16#5bda# => X"0c000028",
		16#5bdb# => X"a86e0000",
		16#5bdc# => X"07ffeca4",
		16#5bdd# => X"a8820000",
		16#5bde# => X"aa0b0000",
		16#5bdf# => X"8562002c",
		16#5be0# => X"bc0b0000",
		16#5be1# => X"10000007",
		16#5be2# => X"a86e0000",
		16#5be3# => X"48005800",
		16#5be4# => X"8482001c",
		16#5be5# => X"bd8b0000",
		16#5be6# => X"10000031",
		16#5be7# => X"15000000",
		16#5be8# => X"9462000c",
		16#5be9# => X"a4630080",
		16#5bea# => X"bc030000",
		16#5beb# => X"0c000028",
		16#5bec# => X"a86e0000",
		16#5bed# => X"84820030",
		16#5bee# => X"bc040000",
		16#5bef# => X"10000009",
		16#5bf0# => X"9c620040",
		16#5bf1# => X"e4041800",
		16#5bf2# => X"10000005",
		16#5bf3# => X"9c600000",
		16#5bf4# => X"07ffeebb",
		16#5bf5# => X"a86e0000",
		16#5bf6# => X"9c600000",
		16#5bf7# => X"d4021830",
		16#5bf8# => X"84820044",
		16#5bf9# => X"bc040000",
		16#5bfa# => X"10000007",
		16#5bfb# => X"9c600000",
		16#5bfc# => X"07ffeeb3",
		16#5bfd# => X"a86e0000",
		16#5bfe# => X"9c600000",
		16#5bff# => X"d4021844",
		16#5c00# => X"9c600000",
		16#5c01# => X"dc02180c",
		16#5c02# => X"07ffee43",
		16#5c03# => X"15000000",
		16#5c04# => X"9c210010",
		16#5c05# => X"a9700000",
		16#5c06# => X"8521fffc",
		16#5c07# => X"8441fff0",
		16#5c08# => X"85c1fff4",
		16#5c09# => X"44004800",
		16#5c0a# => X"8601fff8",
		16#5c0b# => X"07ffed83",
		16#5c0c# => X"a86e0000",
		16#5c0d# => X"9a02000c",
		16#5c0e# => X"bc300000",
		16#5c0f# => X"13ffffcd",
		16#5c10# => X"a86e0000",
		16#5c11# => X"03fffff1",
		16#5c12# => X"15000000",
		16#5c13# => X"07ffee9c",
		16#5c14# => X"84820010",
		16#5c15# => X"03ffffd9",
		16#5c16# => X"84820030",
		16#5c17# => X"03ffffd1",
		16#5c18# => X"9e00ffff",
		16#5c19# => X"a8830000",
		16#5c1a# => X"18600001",
		16#5c1b# => X"d7e14ffc",
		16#5c1c# => X"a863ade4",
		16#5c1d# => X"9c21fffc",
		16#5c1e# => X"84630000",
		16#5c1f# => X"9c210004",
		16#5c20# => X"8521fffc",
		16#5c21# => X"03ffffa4",
		16#5c22# => X"15000000",
		16#5c23# => X"d7e1b7f8",
		16#5c24# => X"aac30000",
		16#5c25# => X"9865000c",
		16#5c26# => X"d7e117e4",
		16#5c27# => X"d7e1a7f4",
		16#5c28# => X"d7e14ffc",
		16#5c29# => X"d7e177e8",
		16#5c2a# => X"d7e187ec",
		16#5c2b# => X"d7e197f0",
		16#5c2c# => X"a8450000",
		16#5c2d# => X"a4a32000",
		16#5c2e# => X"9c21ffe0",
		16#5c2f# => X"bc250000",
		16#5c30# => X"10000007",
		16#5c31# => X"aa840000",
		16#5c32# => X"84820064",
		16#5c33# => X"a8632000",
		16#5c34# => X"a8842000",
		16#5c35# => X"dc02180c",
		16#5c36# => X"d4022064",
		16#5c37# => X"bdb40000",
		16#5c38# => X"1000003e",
		16#5c39# => X"18600001",
		16#5c3a# => X"a863b794",
		16#5c3b# => X"84630000",
		16#5c3c# => X"ac630001",
		16#5c3d# => X"e0801802",
		16#5c3e# => X"e0641804",
		16#5c3f# => X"bd830000",
		16#5c40# => X"10000036",
		16#5c41# => X"bd5400ff",
		16#5c42# => X"10000034",
		16#5c43# => X"9e400001",
		16#5c44# => X"d801a003",
		16#5c45# => X"9dc10003",
		16#5c46# => X"0000000c",
		16#5c47# => X"9e000000",
		16#5c48# => X"8c6e0000",
		16#5c49# => X"84820000",
		16#5c4a# => X"d8041800",
		16#5c4b# => X"84c20000",
		16#5c4c# => X"9cc60001",
		16#5c4d# => X"d4023000",
		16#5c4e# => X"9e100001",
		16#5c4f# => X"e4909000",
		16#5c50# => X"0c000032",
		16#5c51# => X"9dce0001",
		16#5c52# => X"84c20008",
		16#5c53# => X"9cc6ffff",
		16#5c54# => X"bd660000",
		16#5c55# => X"13fffff3",
		16#5c56# => X"d4023008",
		16#5c57# => X"84620018",
		16#5c58# => X"e5861800",
		16#5c59# => X"1000002f",
		16#5c5a# => X"15000000",
		16#5c5b# => X"8c8e0000",
		16#5c5c# => X"84620000",
		16#5c5d# => X"d8032000",
		16#5c5e# => X"84820000",
		16#5c5f# => X"8cc40000",
		16#5c60# => X"ac66ffff",
		16#5c61# => X"9ca40001",
		16#5c62# => X"e0801802",
		16#5c63# => X"bc06000a",
		16#5c64# => X"1000002e",
		16#5c65# => X"e0641804",
		16#5c66# => X"ac63ffff",
		16#5c67# => X"d4022800",
		16#5c68# => X"b8c3005f",
		16#5c69# => X"bc260000",
		16#5c6a# => X"0fffffe5",
		16#5c6b# => X"9e100001",
		16#5c6c# => X"9d60ffff",
		16#5c6d# => X"9c210020",
		16#5c6e# => X"8521fffc",
		16#5c6f# => X"8441ffe4",
		16#5c70# => X"85c1ffe8",
		16#5c71# => X"8601ffec",
		16#5c72# => X"8641fff0",
		16#5c73# => X"8681fff4",
		16#5c74# => X"44004800",
		16#5c75# => X"86c1fff8",
		16#5c76# => X"9dc10003",
		16#5c77# => X"a8760000",
		16#5c78# => X"a88e0000",
		16#5c79# => X"a8b40000",
		16#5c7a# => X"040000af",
		16#5c7b# => X"9cc2005c",
		16#5c7c# => X"bc2bffff",
		16#5c7d# => X"0c000007",
		16#5c7e# => X"aa4b0000",
		16#5c7f# => X"bc2b0000",
		16#5c80# => X"13ffffd2",
		16#5c81# => X"9e000000",
		16#5c82# => X"03ffffeb",
		16#5c83# => X"a9740000",
		16#5c84# => X"9462000c",
		16#5c85# => X"a8630040",
		16#5c86# => X"03ffffe7",
		16#5c87# => X"dc02180c",
		16#5c88# => X"8c8e0000",
		16#5c89# => X"a8760000",
		16#5c8a# => X"07ffe287",
		16#5c8b# => X"a8a20000",
		16#5c8c# => X"ad6bffff",
		16#5c8d# => X"e0c05802",
		16#5c8e# => X"e0c65804",
		16#5c8f# => X"acc6ffff",
		16#5c90# => X"03ffffd9",
		16#5c91# => X"b8c6005f",
		16#5c92# => X"a8760000",
		16#5c93# => X"03fffff7",
		16#5c94# => X"a8860000",
		16#5c95# => X"d7e187f8",
		16#5c96# => X"1a000001",
		16#5c97# => X"d7e117f0",
		16#5c98# => X"aa10ade4",
		16#5c99# => X"d7e177f4",
		16#5c9a# => X"d7e14ffc",
		16#5c9b# => X"a9c30000",
		16#5c9c# => X"84700000",
		16#5c9d# => X"9c21fff0",
		16#5c9e# => X"bc030000",
		16#5c9f# => X"10000009",
		16#5ca0# => X"a8440000",
		16#5ca1# => X"84830038",
		16#5ca2# => X"bc240000",
		16#5ca3# => X"10000005",
		16#5ca4# => X"15000000",
		16#5ca5# => X"07ffece9",
		16#5ca6# => X"15000000",
		16#5ca7# => X"84700000",
		16#5ca8# => X"9c210010",
		16#5ca9# => X"a88e0000",
		16#5caa# => X"a8a20000",
		16#5cab# => X"8521fffc",
		16#5cac# => X"8441fff0",
		16#5cad# => X"85c1fff4",
		16#5cae# => X"03ffff75",
		16#5caf# => X"8601fff8",
		16#5cb0# => X"d7e117f4",
		16#5cb1# => X"18400001",
		16#5cb2# => X"d7e177f8",
		16#5cb3# => X"a842c508",
		16#5cb4# => X"a9c30000",
		16#5cb5# => X"a8640000",
		16#5cb6# => X"a8850000",
		16#5cb7# => X"9ca00000",
		16#5cb8# => X"d7e14ffc",
		16#5cb9# => X"d4022800",
		16#5cba# => X"0400010b",
		16#5cbb# => X"9c21fff4",
		16#5cbc# => X"bc2bffff",
		16#5cbd# => X"0c000007",
		16#5cbe# => X"15000000",
		16#5cbf# => X"9c21000c",
		16#5cc0# => X"8521fffc",
		16#5cc1# => X"8441fff4",
		16#5cc2# => X"44004800",
		16#5cc3# => X"85c1fff8",
		16#5cc4# => X"84420000",
		16#5cc5# => X"bc020000",
		16#5cc6# => X"13fffff9",
		16#5cc7# => X"15000000",
		16#5cc8# => X"d40e1000",
		16#5cc9# => X"9c21000c",
		16#5cca# => X"8521fffc",
		16#5ccb# => X"8441fff4",
		16#5ccc# => X"44004800",
		16#5ccd# => X"85c1fff8",
		16#5cce# => X"d7e117f4",
		16#5ccf# => X"18400001",
		16#5cd0# => X"d7e177f8",
		16#5cd1# => X"a842c508",
		16#5cd2# => X"a9c30000",
		16#5cd3# => X"a8640000",
		16#5cd4# => X"9c800000",
		16#5cd5# => X"d7e14ffc",
		16#5cd6# => X"d4022000",
		16#5cd7# => X"04000179",
		16#5cd8# => X"9c21fff4",
		16#5cd9# => X"bc2bffff",
		16#5cda# => X"0c000007",
		16#5cdb# => X"15000000",
		16#5cdc# => X"9c21000c",
		16#5cdd# => X"8521fffc",
		16#5cde# => X"8441fff4",
		16#5cdf# => X"44004800",
		16#5ce0# => X"85c1fff8",
		16#5ce1# => X"84420000",
		16#5ce2# => X"bc020000",
		16#5ce3# => X"13fffff9",
		16#5ce4# => X"15000000",
		16#5ce5# => X"d40e1000",
		16#5ce6# => X"9c21000c",
		16#5ce7# => X"8521fffc",
		16#5ce8# => X"8441fff4",
		16#5ce9# => X"44004800",
		16#5cea# => X"85c1fff8",
		16#5ceb# => X"d7e117f4",
		16#5cec# => X"18400001",
		16#5ced# => X"d7e177f8",
		16#5cee# => X"a842c508",
		16#5cef# => X"a9c30000",
		16#5cf0# => X"a8640000",
		16#5cf1# => X"a8850000",
		16#5cf2# => X"a8a60000",
		16#5cf3# => X"9cc00000",
		16#5cf4# => X"d7e14ffc",
		16#5cf5# => X"d4023000",
		16#5cf6# => X"04000183",
		16#5cf7# => X"9c21fff4",
		16#5cf8# => X"bc2bffff",
		16#5cf9# => X"0c000007",
		16#5cfa# => X"15000000",
		16#5cfb# => X"9c21000c",
		16#5cfc# => X"8521fffc",
		16#5cfd# => X"8441fff4",
		16#5cfe# => X"44004800",
		16#5cff# => X"85c1fff8",
		16#5d00# => X"84420000",
		16#5d01# => X"bc020000",
		16#5d02# => X"13fffff9",
		16#5d03# => X"15000000",
		16#5d04# => X"d40e1000",
		16#5d05# => X"9c21000c",
		16#5d06# => X"8521fffc",
		16#5d07# => X"8441fff4",
		16#5d08# => X"44004800",
		16#5d09# => X"85c1fff8",
		16#5d0a# => X"d7e117f4",
		16#5d0b# => X"18400001",
		16#5d0c# => X"d7e177f8",
		16#5d0d# => X"a842c508",
		16#5d0e# => X"a9c30000",
		16#5d0f# => X"a8640000",
		16#5d10# => X"a8850000",
		16#5d11# => X"a8a60000",
		16#5d12# => X"9cc00000",
		16#5d13# => X"d7e14ffc",
		16#5d14# => X"d4023000",
		16#5d15# => X"04000186",
		16#5d16# => X"9c21fff4",
		16#5d17# => X"bc2bffff",
		16#5d18# => X"0c000007",
		16#5d19# => X"15000000",
		16#5d1a# => X"9c21000c",
		16#5d1b# => X"8521fffc",
		16#5d1c# => X"8441fff4",
		16#5d1d# => X"44004800",
		16#5d1e# => X"85c1fff8",
		16#5d1f# => X"84420000",
		16#5d20# => X"bc020000",
		16#5d21# => X"13fffff9",
		16#5d22# => X"15000000",
		16#5d23# => X"d40e1000",
		16#5d24# => X"9c21000c",
		16#5d25# => X"8521fffc",
		16#5d26# => X"8441fff4",
		16#5d27# => X"44004800",
		16#5d28# => X"85c1fff8",
		16#5d29# => X"d7e117e8",
		16#5d2a# => X"d7e177ec",
		16#5d2b# => X"d7e187f0",
		16#5d2c# => X"d7e197f4",
		16#5d2d# => X"d7e14ffc",
		16#5d2e# => X"d7e1a7f8",
		16#5d2f# => X"a8440000",
		16#5d30# => X"9c21ffdc",
		16#5d31# => X"aa030000",
		16#5d32# => X"a9c50000",
		16#5d33# => X"bc240000",
		16#5d34# => X"0c00001a",
		16#5d35# => X"aa460000",
		16#5d36# => X"18600001",
		16#5d37# => X"a863b7d8",
		16#5d38# => X"07fff040",
		16#5d39# => X"86830000",
		16#5d3a# => X"a8700000",
		16#5d3b# => X"a8820000",
		16#5d3c# => X"a8ae0000",
		16#5d3d# => X"a8cb0000",
		16#5d3e# => X"4800a000",
		16#5d3f# => X"a8f20000",
		16#5d40# => X"bc2bffff",
		16#5d41# => X"10000005",
		16#5d42# => X"9c400000",
		16#5d43# => X"d4121000",
		16#5d44# => X"9c40008a",
		16#5d45# => X"d4101000",
		16#5d46# => X"9c210024",
		16#5d47# => X"8521fffc",
		16#5d48# => X"8441ffe8",
		16#5d49# => X"85c1ffec",
		16#5d4a# => X"8601fff0",
		16#5d4b# => X"8641fff4",
		16#5d4c# => X"44004800",
		16#5d4d# => X"8681fff8",
		16#5d4e# => X"18600001",
		16#5d4f# => X"a863b7d8",
		16#5d50# => X"07fff028",
		16#5d51# => X"85c30000",
		16#5d52# => X"a8700000",
		16#5d53# => X"a8810000",
		16#5d54# => X"a8a20000",
		16#5d55# => X"a8cb0000",
		16#5d56# => X"48007000",
		16#5d57# => X"a8f20000",
		16#5d58# => X"03ffffe9",
		16#5d59# => X"bc2bffff",
		16#5d5a# => X"d7e117e4",
		16#5d5b# => X"d7e177e8",
		16#5d5c# => X"d7e197f0",
		16#5d5d# => X"d7e14ffc",
		16#5d5e# => X"d7e187ec",
		16#5d5f# => X"d7e1a7f4",
		16#5d60# => X"d7e1b7f8",
		16#5d61# => X"a8430000",
		16#5d62# => X"9c21ffd8",
		16#5d63# => X"aa440000",
		16#5d64# => X"bc230000",
		16#5d65# => X"0c00001f",
		16#5d66# => X"a9c50000",
		16#5d67# => X"1a000001",
		16#5d68# => X"18600001",
		16#5d69# => X"aa10ade4",
		16#5d6a# => X"a863b7d8",
		16#5d6b# => X"86d00000",
		16#5d6c# => X"07fff00c",
		16#5d6d# => X"86830000",
		16#5d6e# => X"a8760000",
		16#5d6f# => X"a8820000",
		16#5d70# => X"a8b20000",
		16#5d71# => X"a8cb0000",
		16#5d72# => X"4800a000",
		16#5d73# => X"a8ee0000",
		16#5d74# => X"bc2bffff",
		16#5d75# => X"10000006",
		16#5d76# => X"9c600000",
		16#5d77# => X"84500000",
		16#5d78# => X"d40e1800",
		16#5d79# => X"9c60008a",
		16#5d7a# => X"d4021800",
		16#5d7b# => X"9c210028",
		16#5d7c# => X"8521fffc",
		16#5d7d# => X"8441ffe4",
		16#5d7e# => X"85c1ffe8",
		16#5d7f# => X"8601ffec",
		16#5d80# => X"8641fff0",
		16#5d81# => X"8681fff4",
		16#5d82# => X"44004800",
		16#5d83# => X"86c1fff8",
		16#5d84# => X"1a000001",
		16#5d85# => X"18600001",
		16#5d86# => X"aa10ade4",
		16#5d87# => X"a863b7d8",
		16#5d88# => X"86900000",
		16#5d89# => X"07ffefef",
		16#5d8a# => X"86430000",
		16#5d8b# => X"a8740000",
		16#5d8c# => X"a8810000",
		16#5d8d# => X"a8a20000",
		16#5d8e# => X"a8cb0000",
		16#5d8f# => X"48009000",
		16#5d90# => X"a8ee0000",
		16#5d91# => X"03ffffe4",
		16#5d92# => X"bc2bffff",
		16#5d93# => X"bc040000",
		16#5d94# => X"10000006",
		16#5d95# => X"bca500ff",
		16#5d96# => X"0c000006",
		16#5d97# => X"15000000",
		16#5d98# => X"d8042800",
		16#5d99# => X"9c800001",
		16#5d9a# => X"44004800",
		16#5d9b# => X"a9640000",
		16#5d9c# => X"9ca0008a",
		16#5d9d# => X"9c80ffff",
		16#5d9e# => X"03fffffc",
		16#5d9f# => X"d4032800",
		16#5da0# => X"d7e187f0",
		16#5da1# => X"aa030000",
		16#5da2# => X"18600001",
		16#5da3# => X"d7e14ffc",
		16#5da4# => X"d7e117e8",
		16#5da5# => X"d7e177ec",
		16#5da6# => X"d7e197f4",
		16#5da7# => X"d7e1a7f8",
		16#5da8# => X"a863b7d8",
		16#5da9# => X"9c21ffe8",
		16#5daa# => X"aa860000",
		16#5dab# => X"a9c40000",
		16#5dac# => X"a8450000",
		16#5dad# => X"07ffefcb",
		16#5dae# => X"86430000",
		16#5daf# => X"9c210018",
		16#5db0# => X"a8700000",
		16#5db1# => X"a88e0000",
		16#5db2# => X"a8a20000",
		16#5db3# => X"a8f40000",
		16#5db4# => X"a8cb0000",
		16#5db5# => X"8521fffc",
		16#5db6# => X"8441ffe8",
		16#5db7# => X"85c1ffec",
		16#5db8# => X"8601fff0",
		16#5db9# => X"8681fff8",
		16#5dba# => X"44009000",
		16#5dbb# => X"8641fff4",
		16#5dbc# => X"15000001",
		16#5dbd# => X"00000000",
		16#5dbe# => X"15000000",
		16#5dbf# => X"18600001",
		16#5dc0# => X"9c800009",
		16#5dc1# => X"a863c508",
		16#5dc2# => X"9d60ffff",
		16#5dc3# => X"44004800",
		16#5dc4# => X"d4032000",
		16#5dc5# => X"e0a01802",
		16#5dc6# => X"e0a51804",
		16#5dc7# => X"bd850000",
		16#5dc8# => X"0c00000c",
		16#5dc9# => X"18a00001",
		16#5dca# => X"aca30001",
		16#5dcb# => X"e0c02802",
		16#5dcc# => X"e0a62804",
		16#5dcd# => X"bd650000",
		16#5dce# => X"0c00000f",
		16#5dcf# => X"ac630002",
		16#5dd0# => X"9c602000",
		16#5dd1# => X"9d600000",
		16#5dd2# => X"44004800",
		16#5dd3# => X"d4041804",
		16#5dd4# => X"a8a57da8",
		16#5dd5# => X"84a50000",
		16#5dd6# => X"e0c02802",
		16#5dd7# => X"e0a62804",
		16#5dd8# => X"bd850000",
		16#5dd9# => X"0ffffff2",
		16#5dda# => X"aca30001",
		16#5ddb# => X"03fffff6",
		16#5ddc# => X"9c602000",
		16#5ddd# => X"e0a01802",
		16#5dde# => X"e0651804",
		16#5ddf# => X"bd830000",
		16#5de0# => X"0ffffff1",
		16#5de1# => X"9c602000",
		16#5de2# => X"18600001",
		16#5de3# => X"9c800009",
		16#5de4# => X"a863c508",
		16#5de5# => X"9d60ffff",
		16#5de6# => X"44004800",
		16#5de7# => X"d4032000",
		16#5de8# => X"19000001",
		16#5de9# => X"9c800000",
		16#5dea# => X"a908ade4",
		16#5deb# => X"d7e14ffc",
		16#5dec# => X"84a80000",
		16#5ded# => X"d7e117f8",
		16#5dee# => X"9ce50014",
		16#5def# => X"9da502ec",
		16#5df0# => X"d8072018",
		16#5df1# => X"9d850354",
		16#5df2# => X"9d6503bc",
		16#5df3# => X"84680000",
		16#5df4# => X"d4056804",
		16#5df5# => X"d4052000",
		16#5df6# => X"d4056008",
		16#5df7# => X"d405580c",
		16#5df8# => X"d4052010",
		16#5df9# => X"18a00001",
		16#5dfa# => X"9cc3007c",
		16#5dfb# => X"a8a58894",
		16#5dfc# => X"d4032030",
		16#5dfd# => X"d4032834",
		16#5dfe# => X"d4032038",
		16#5dff# => X"d403203c",
		16#5e00# => X"d4032040",
		16#5e01# => X"d4032044",
		16#5e02# => X"d4032048",
		16#5e03# => X"d403204c",
		16#5e04# => X"d4032050",
		16#5e05# => X"d4032054",
		16#5e06# => X"d4032058",
		16#5e07# => X"d403205c",
		16#5e08# => X"d8032060",
		16#5e09# => X"d4072000",
		16#5e0a# => X"d4072004",
		16#5e0b# => X"d4072008",
		16#5e0c# => X"d407200c",
		16#5e0d# => X"d4072010",
		16#5e0e# => X"d4072014",
		16#5e0f# => X"d4062000",
		16#5e10# => X"d4062004",
		16#5e11# => X"d4062008",
		16#5e12# => X"d406200c",
		16#5e13# => X"d4062010",
		16#5e14# => X"9c400000",
		16#5e15# => X"84a80000",
		16#5e16# => X"9c600001",
		16#5e17# => X"d40520a0",
		16#5e18# => X"d40510a4",
		16#5e19# => X"d40518a8",
		16#5e1a# => X"9c60330e",
		16#5e1b# => X"9c40abcd",
		16#5e1c# => X"dc0518ac",
		16#5e1d# => X"9c601234",
		16#5e1e# => X"dc0510ae",
		16#5e1f# => X"dc0518b0",
		16#5e20# => X"9c40e66d",
		16#5e21# => X"9c60deec",
		16#5e22# => X"dc0510b2",
		16#5e23# => X"dc0518b4",
		16#5e24# => X"9c400005",
		16#5e25# => X"9c60000b",
		16#5e26# => X"dc0510b6",
		16#5e27# => X"dc0518b8",
		16#5e28# => X"d40520bc",
		16#5e29# => X"d40520c0",
		16#5e2a# => X"d40520c4",
		16#5e2b# => X"d40520c8",
		16#5e2c# => X"d40520cc",
		16#5e2d# => X"d40520d0",
		16#5e2e# => X"d40520f8",
		16#5e2f# => X"d40520fc",
		16#5e30# => X"d4052100",
		16#5e31# => X"d4052104",
		16#5e32# => X"d4052108",
		16#5e33# => X"d405210c",
		16#5e34# => X"d4052110",
		16#5e35# => X"d4052114",
		16#5e36# => X"d4052118",
		16#5e37# => X"d405211c",
		16#5e38# => X"d80520d4",
		16#5e39# => X"d80520dc",
		16#5e3a# => X"d40520f4",
		16#5e3b# => X"9c21fff8",
		16#5e3c# => X"d4062014",
		16#5e3d# => X"d4062018",
		16#5e3e# => X"d406201c",
		16#5e3f# => X"d4062020",
		16#5e40# => X"d4052148",
		16#5e41# => X"d405214c",
		16#5e42# => X"d4052150",
		16#5e43# => X"d4052154",
		16#5e44# => X"d40522d4",
		16#5e45# => X"d40521d4",
		16#5e46# => X"d40522dc",
		16#5e47# => X"d40522e0",
		16#5e48# => X"d40522e4",
		16#5e49# => X"d40522e8",
		16#5e4a# => X"9c210008",
		16#5e4b# => X"9c6502ec",
		16#5e4c# => X"8521fffc",
		16#5e4d# => X"9ca00138",
		16#5e4e# => X"03fff0ab",
		16#5e4f# => X"8441fff8",
		16#5e50# => X"e0801802",
		16#5e51# => X"d7e14ffc",
		16#5e52# => X"e0841804",
		16#5e53# => X"bd840000",
		16#5e54# => X"0c00000d",
		16#5e55# => X"9c21fffc",
		16#5e56# => X"ac830002",
		16#5e57# => X"e0a02002",
		16#5e58# => X"e0852004",
		16#5e59# => X"bd640000",
		16#5e5a# => X"0c000013",
		16#5e5b# => X"15000000",
		16#5e5c# => X"9c800001",
		16#5e5d# => X"9c210004",
		16#5e5e# => X"8521fffc",
		16#5e5f# => X"44004800",
		16#5e60# => X"a9640000",
		16#5e61# => X"18a00001",
		16#5e62# => X"a8a57da8",
		16#5e63# => X"84a50000",
		16#5e64# => X"e0c02802",
		16#5e65# => X"e0a62804",
		16#5e66# => X"bd850000",
		16#5e67# => X"0fffffef",
		16#5e68# => X"9c800001",
		16#5e69# => X"9c210004",
		16#5e6a# => X"8521fffc",
		16#5e6b# => X"44004800",
		16#5e6c# => X"a9640000",
		16#5e6d# => X"ac630001",
		16#5e6e# => X"e0801802",
		16#5e6f# => X"e0641804",
		16#5e70# => X"bd630000",
		16#5e71# => X"13ffffeb",
		16#5e72# => X"15000000",
		16#5e73# => X"040000f9",
		16#5e74# => X"15000000",
		16#5e75# => X"9c600009",
		16#5e76# => X"9c80ffff",
		16#5e77# => X"03ffffe6",
		16#5e78# => X"d40b1800",
		16#5e79# => X"e0801802",
		16#5e7a# => X"e0841804",
		16#5e7b# => X"bd840000",
		16#5e7c# => X"0c00000a",
		16#5e7d# => X"18800001",
		16#5e7e# => X"ac830002",
		16#5e7f# => X"e0a02002",
		16#5e80# => X"e0852004",
		16#5e81# => X"bd640000",
		16#5e82# => X"0c00000e",
		16#5e83# => X"15000000",
		16#5e84# => X"44004800",
		16#5e85# => X"9d600000",
		16#5e86# => X"9d600000",
		16#5e87# => X"a8847da8",
		16#5e88# => X"84840000",
		16#5e89# => X"e0a02002",
		16#5e8a# => X"e0852004",
		16#5e8b# => X"e5845800",
		16#5e8c# => X"0ffffff2",
		16#5e8d# => X"15000000",
		16#5e8e# => X"44004800",
		16#5e8f# => X"15000000",
		16#5e90# => X"ac630001",
		16#5e91# => X"e0801802",
		16#5e92# => X"e0641804",
		16#5e93# => X"bd630000",
		16#5e94# => X"13fffff0",
		16#5e95# => X"9c800009",
		16#5e96# => X"18600001",
		16#5e97# => X"a863c508",
		16#5e98# => X"9d60ffff",
		16#5e99# => X"44004800",
		16#5e9a# => X"d4032000",
		16#5e9b# => X"d7e177f4",
		16#5e9c# => X"d7e187f8",
		16#5e9d# => X"d7e14ffc",
		16#5e9e# => X"d7e117f0",
		16#5e9f# => X"aa040000",
		16#5ea0# => X"9c21fff0",
		16#5ea1# => X"bc230000",
		16#5ea2# => X"1000001f",
		16#5ea3# => X"a9c50000",
		16#5ea4# => X"18400001",
		16#5ea5# => X"a8427da8",
		16#5ea6# => X"84420000",
		16#5ea7# => X"bc020000",
		16#5ea8# => X"10000012",
		16#5ea9# => X"bda50000",
		16#5eaa# => X"0c000008",
		16#5eab# => X"a8430000",
		16#5eac# => X"0000000f",
		16#5ead# => X"9c210010",
		16#5eae# => X"9c420001",
		16#5eaf# => X"e54e1000",
		16#5eb0# => X"0c00000a",
		16#5eb1# => X"15000000",
		16#5eb2# => X"04000073",
		16#5eb3# => X"15000000",
		16#5eb4# => X"b96b0018",
		16#5eb5# => X"e0701000",
		16#5eb6# => X"b96b0098",
		16#5eb7# => X"bc0b000a",
		16#5eb8# => X"0ffffff6",
		16#5eb9# => X"d8035800",
		16#5eba# => X"9c210010",
		16#5ebb# => X"a9620000",
		16#5ebc# => X"8521fffc",
		16#5ebd# => X"8441fff0",
		16#5ebe# => X"85c1fff4",
		16#5ebf# => X"44004800",
		16#5ec0# => X"8601fff8",
		16#5ec1# => X"18600001",
		16#5ec2# => X"9c800009",
		16#5ec3# => X"a863c508",
		16#5ec4# => X"9c40ffff",
		16#5ec5# => X"03fffff5",
		16#5ec6# => X"d4032000",
		16#5ec7# => X"18800001",
		16#5ec8# => X"18a00001",
		16#5ec9# => X"a884b7dc",
		16#5eca# => X"a8a5adc4",
		16#5ecb# => X"85640000",
		16#5ecc# => X"84a50000",
		16#5ecd# => X"e06b1800",
		16#5ece# => X"d7e117fc",
		16#5ecf# => X"e0a51802",
		16#5ed0# => X"18400001",
		16#5ed1# => X"e5a51000",
		16#5ed2# => X"0c00000a",
		16#5ed3# => X"9c21fffc",
		16#5ed4# => X"18600001",
		16#5ed5# => X"9c80000c",
		16#5ed6# => X"a863c508",
		16#5ed7# => X"9d60ffff",
		16#5ed8# => X"d4032000",
		16#5ed9# => X"9c210004",
		16#5eda# => X"44004800",
		16#5edb# => X"8441fffc",
		16#5edc# => X"d4041800",
		16#5edd# => X"9c210004",
		16#5ede# => X"44004800",
		16#5edf# => X"8441fffc",
		16#5ee0# => X"d7e117f8",
		16#5ee1# => X"18400001",
		16#5ee2# => X"9c80ffc7",
		16#5ee3# => X"a8427da8",
		16#5ee4# => X"d7e14ffc",
		16#5ee5# => X"84620000",
		16#5ee6# => X"9c21fff8",
		16#5ee7# => X"9c630002",
		16#5ee8# => X"d8032000",
		16#5ee9# => X"9c800000",
		16#5eea# => X"84620000",
		16#5eeb# => X"9c630001",
		16#5eec# => X"d8032000",
		16#5eed# => X"9c800003",
		16#5eee# => X"84620000",
		16#5eef# => X"9c630003",
		16#5ef0# => X"d8032000",
		16#5ef1# => X"18600001",
		16#5ef2# => X"18800001",
		16#5ef3# => X"a8637da4",
		16#5ef4# => X"a8847dac",
		16#5ef5# => X"84630000",
		16#5ef6# => X"07ffc6d6",
		16#5ef7# => X"84840000",
		16#5ef8# => X"84620000",
		16#5ef9# => X"9d6b0008",
		16#5efa# => X"9c630003",
		16#5efb# => X"b96b0044",
		16#5efc# => X"8ca30000",
		16#5efd# => X"a8a50080",
		16#5efe# => X"a48b00ff",
		16#5eff# => X"d8032800",
		16#5f00# => X"b96b0088",
		16#5f01# => X"84620000",
		16#5f02# => X"d8032000",
		16#5f03# => X"a56b00ff",
		16#5f04# => X"84620000",
		16#5f05# => X"9c630001",
		16#5f06# => X"d8035800",
		16#5f07# => X"84420000",
		16#5f08# => X"9c420003",
		16#5f09# => X"8c620000",
		16#5f0a# => X"a463007f",
		16#5f0b# => X"d8021800",
		16#5f0c# => X"9c210008",
		16#5f0d# => X"8521fffc",
		16#5f0e# => X"44004800",
		16#5f0f# => X"8441fff8",
		16#5f10# => X"18a00001",
		16#5f11# => X"b8630018",
		16#5f12# => X"a8a57da8",
		16#5f13# => X"84c50000",
		16#5f14# => X"b8e30098",
		16#5f15# => X"9c860005",
		16#5f16# => X"8c640000",
		16#5f17# => X"a4630020",
		16#5f18# => X"bc030000",
		16#5f19# => X"13fffffd",
		16#5f1a# => X"a46700ff",
		16#5f1b# => X"d8061800",
		16#5f1c# => X"84850000",
		16#5f1d# => X"9c840005",
		16#5f1e# => X"8c640000",
		16#5f1f# => X"a4630060",
		16#5f20# => X"bc230060",
		16#5f21# => X"13fffffd",
		16#5f22# => X"15000000",
		16#5f23# => X"44004800",
		16#5f24# => X"15000000",
		16#5f25# => X"18600001",
		16#5f26# => X"a8637da8",
		16#5f27# => X"84a30000",
		16#5f28# => X"9c850005",
		16#5f29# => X"8c640000",
		16#5f2a# => X"a4630001",
		16#5f2b# => X"bc030000",
		16#5f2c# => X"13fffffd",
		16#5f2d# => X"15000000",
		16#5f2e# => X"8d650000",
		16#5f2f# => X"b96b0018",
		16#5f30# => X"44004800",
		16#5f31# => X"b96b0098",
		16#5f32# => X"d7e187f4",
		16#5f33# => X"d7e197f8",
		16#5f34# => X"d7e14ffc",
		16#5f35# => X"d7e117ec",
		16#5f36# => X"d7e177f0",
		16#5f37# => X"9c63ffff",
		16#5f38# => X"9c21ffec",
		16#5f39# => X"aa440000",
		16#5f3a# => X"bc430001",
		16#5f3b# => X"1000001f",
		16#5f3c# => X"aa050000",
		16#5f3d# => X"bd450000",
		16#5f3e# => X"0c000014",
		16#5f3f# => X"19c00001",
		16#5f40# => X"9c400000",
		16#5f41# => X"00000007",
		16#5f42# => X"a9ce7da8",
		16#5f43# => X"15000004",
		16#5f44# => X"9c420001",
		16#5f45# => X"e5501000",
		16#5f46# => X"0c00000c",
		16#5f47# => X"15000000",
		16#5f48# => X"848e0000",
		16#5f49# => X"e0721000",
		16#5f4a# => X"bc040000",
		16#5f4b# => X"13fffff8",
		16#5f4c# => X"90630000",
		16#5f4d# => X"07ffffc3",
		16#5f4e# => X"9c420001",
		16#5f4f# => X"e5501000",
		16#5f50# => X"13fffff8",
		16#5f51# => X"15000000",
		16#5f52# => X"9c210014",
		16#5f53# => X"a9700000",
		16#5f54# => X"8521fffc",
		16#5f55# => X"8441ffec",
		16#5f56# => X"85c1fff0",
		16#5f57# => X"8601fff4",
		16#5f58# => X"44004800",
		16#5f59# => X"8641fff8",
		16#5f5a# => X"18400001",
		16#5f5b# => X"9c600009",
		16#5f5c# => X"a842c508",
		16#5f5d# => X"9e00ffff",
		16#5f5e# => X"d4021800",
		16#5f5f# => X"9c210014",
		16#5f60# => X"a9700000",
		16#5f61# => X"8521fffc",
		16#5f62# => X"8441ffec",
		16#5f63# => X"85c1fff0",
		16#5f64# => X"8601fff4",
		16#5f65# => X"44004800",
		16#5f66# => X"8641fff8",
		16#5f67# => X"00000000",
		16#5f68# => X"10000000",
		16#5f69# => X"017d7840",
		16#5f6a# => X"90000000",
		16#5f6b# => X"0001c200",
		16#5f6c# => X"18600001",
		16#5f6d# => X"a863ade4",
		16#5f6e# => X"44004800",
		16#5f6f# => X"85630000",
		16#5f70# => X"9c21fffc",
		16#5f71# => X"d4014800",
		16#5f72# => X"07ffc65a",
		16#5f73# => X"15000000",
		16#5f74# => X"9d670000",
		16#5f75# => X"85210000",
		16#5f76# => X"44004800",
		16#5f77# => X"9c210004",
		16#5f78# => X"9c21fff8",
		16#5f79# => X"d4014800",
		16#5f7a# => X"d4017004",
		16#5f7b# => X"9dc00000",
		16#5f7c# => X"e5830000",
		16#5f7d# => X"0c000004",
		16#5f7e# => X"15000000",
		16#5f7f# => X"9dc00001",
		16#5f80# => X"e0601802",
		16#5f81# => X"e5840000",
		16#5f82# => X"0c000003",
		16#5f83# => X"15000000",
		16#5f84# => X"e0802002",
		16#5f85# => X"07ffc647",
		16#5f86# => X"15000000",
		16#5f87# => X"bc0e0001",
		16#5f88# => X"0c000003",
		16#5f89# => X"9d670000",
		16#5f8a# => X"e1605802",
		16#5f8b# => X"85210000",
		16#5f8c# => X"85c10004",
		16#5f8d# => X"44004800",
		16#5f8e# => X"9c210008",
		16#5f8f# => X"d7e117f8",
		16#5f90# => X"18400001",
		16#5f91# => X"d7e14ffc",
		16#5f92# => X"a842adb4",
		16#5f93# => X"8462fffc",
		16#5f94# => X"bc03ffff",
		16#5f95# => X"10000009",
		16#5f96# => X"9c21fff8",
		16#5f97# => X"9c42fffc",
		16#5f98# => X"48001800",
		16#5f99# => X"9c42fffc",
		16#5f9a# => X"84620000",
		16#5f9b# => X"bc23ffff",
		16#5f9c# => X"13fffffc",
		16#5f9d# => X"15000000",
		16#5f9e# => X"9c210008",
		16#5f9f# => X"8521fffc",
		16#5fa0# => X"44004800",
		16#5fa1# => X"8441fff8",
		16#5fa2# => X"d7e14ffc",
		16#5fa3# => X"9c21fffc",
		16#5fa4# => X"9c210004",
		16#5fa5# => X"8521fffc",
		16#5fa6# => X"44004800",
		16#5fa7# => X"15000000",
		16#5fa8# => X"9c21fffc",
		16#5fa9# => X"d4014800",
		16#5faa# => X"07ffa88f",
		16#5fab# => X"15000000",
		16#5fac# => X"85210000",
		16#5fad# => X"44004800",
		16#5fae# => X"9c210004",
		16#5faf# => X"43505520",
		16#5fb0# => X"25643a20",
		16#5fb1# => X"00366b20",
		16#5fb2# => X"70657266",
		16#5fb3# => X"6f726d61",
		16#5fb4# => X"6e636520",
		16#5fb5# => X"72756e20",
		16#5fb6# => X"70617261",
		16#5fb7# => X"6d657465",
		16#5fb8# => X"72732066",
		16#5fb9# => X"6f722063",
		16#5fba# => X"6f72656d",
		16#5fbb# => X"61726b2e",
		16#5fbc# => X"00366b20",
		16#5fbd# => X"76616c69",
		16#5fbe# => X"64617469",
		16#5fbf# => X"6f6e2072",
		16#5fc0# => X"756e2070",
		16#5fc1# => X"6172616d",
		16#5fc2# => X"65746572",
		16#5fc3# => X"7320666f",
		16#5fc4# => X"7220636f",
		16#5fc5# => X"72656d61",
		16#5fc6# => X"726b2e00",
		16#5fc7# => X"50726f66",
		16#5fc8# => X"696c6520",
		16#5fc9# => X"67656e65",
		16#5fca# => X"72617469",
		16#5fcb# => X"6f6e2072",
		16#5fcc# => X"756e2070",
		16#5fcd# => X"6172616d",
		16#5fce# => X"65746572",
		16#5fcf# => X"7320666f",
		16#5fd0# => X"7220636f",
		16#5fd1# => X"72656d61",
		16#5fd2# => X"726b2e00",
		16#5fd3# => X"324b2070",
		16#5fd4# => X"6572666f",
		16#5fd5# => X"726d616e",
		16#5fd6# => X"63652072",
		16#5fd7# => X"756e2070",
		16#5fd8# => X"6172616d",
		16#5fd9# => X"65746572",
		16#5fda# => X"7320666f",
		16#5fdb# => X"7220636f",
		16#5fdc# => X"72656d61",
		16#5fdd# => X"726b2e00",
		16#5fde# => X"324b2076",
		16#5fdf# => X"616c6964",
		16#5fe0# => X"6174696f",
		16#5fe1# => X"6e207275",
		16#5fe2# => X"6e207061",
		16#5fe3# => X"72616d65",
		16#5fe4# => X"74657273",
		16#5fe5# => X"20666f72",
		16#5fe6# => X"20636f72",
		16#5fe7# => X"656d6172",
		16#5fe8# => X"6b2e005b",
		16#5fe9# => X"25755d45",
		16#5fea# => X"52524f52",
		16#5feb# => X"21206c69",
		16#5fec# => X"73742063",
		16#5fed# => X"72632030",
		16#5fee# => X"78253034",
		16#5fef# => X"78202d20",
		16#5ff0# => X"73686f75",
		16#5ff1# => X"6c642062",
		16#5ff2# => X"65203078",
		16#5ff3# => X"25303478",
		16#5ff4# => X"0a005b25",
		16#5ff5# => X"755d4552",
		16#5ff6# => X"524f5221",
		16#5ff7# => X"206d6174",
		16#5ff8# => X"72697820",
		16#5ff9# => X"63726320",
		16#5ffa# => X"30782530",
		16#5ffb# => X"3478202d",
		16#5ffc# => X"2073686f",
		16#5ffd# => X"756c6420",
		16#5ffe# => X"62652030",
		16#5fff# => X"78253034",
		16#6000# => X"780a005b",
		16#6001# => X"25755d45",
		16#6002# => X"52524f52",
		16#6003# => X"21207374",
		16#6004# => X"61746520",
		16#6005# => X"63726320",
		16#6006# => X"30782530",
		16#6007# => X"3478202d",
		16#6008# => X"2073686f",
		16#6009# => X"756c6420",
		16#600a# => X"62652030",
		16#600b# => X"78253034",
		16#600c# => X"780a0043",
		16#600d# => X"6f72654d",
		16#600e# => X"61726b20",
		16#600f# => X"53697a65",
		16#6010# => X"20202020",
		16#6011# => X"3a20256c",
		16#6012# => X"750a0054",
		16#6013# => X"6f74616c",
		16#6014# => X"20746963",
		16#6015# => X"6b732020",
		16#6016# => X"20202020",
		16#6017# => X"3a20256c",
		16#6018# => X"750a0054",
		16#6019# => X"6f74616c",
		16#601a# => X"2074696d",
		16#601b# => X"65202873",
		16#601c# => X"65637329",
		16#601d# => X"3a202566",
		16#601e# => X"0a004974",
		16#601f# => X"65726174",
		16#6020# => X"696f6e73",
		16#6021# => X"2f536563",
		16#6022# => X"2020203a",
		16#6023# => X"2025660a",
		16#6024# => X"00455252",
		16#6025# => X"4f522120",
		16#6026# => X"4d757374",
		16#6027# => X"20657865",
		16#6028# => X"63757465",
		16#6029# => X"20666f72",
		16#602a# => X"20617420",
		16#602b# => X"6c656173",
		16#602c# => X"74203130",
		16#602d# => X"20736563",
		16#602e# => X"7320666f",
		16#602f# => X"72206120",
		16#6030# => X"76616c69",
		16#6031# => X"64207265",
		16#6032# => X"73756c74",
		16#6033# => X"21004974",
		16#6034# => X"65726174",
		16#6035# => X"696f6e73",
		16#6036# => X"20202020",
		16#6037# => X"2020203a",
		16#6038# => X"20256c75",
		16#6039# => X"0a00436f",
		16#603a# => X"6d70696c",
		16#603b# => X"65722076",
		16#603c# => X"65727369",
		16#603d# => X"6f6e203a",
		16#603e# => X"2025730a",
		16#603f# => X"00474343",
		16#6040# => X"342e352e",
		16#6041# => X"312d6f72",
		16#6042# => X"33322d31",
		16#6043# => X"2e307263",
		16#6044# => X"3400436f",
		16#6045# => X"6d70696c",
		16#6046# => X"65722066",
		16#6047# => X"6c616773",
		16#6048# => X"2020203a",
		16#6049# => X"2025730a",
		16#604a# => X"002d4f33",
		16#604b# => X"202d6d68",
		16#604c# => X"6172642d",
		16#604d# => X"6d756c20",
		16#604e# => X"2d6d736f",
		16#604f# => X"66742d64",
		16#6050# => X"6976202d",
		16#6051# => X"6d736f66",
		16#6052# => X"742d666c",
		16#6053# => X"6f617420",
		16#6054# => X"2d445553",
		16#6055# => X"455f504e",
		16#6056# => X"54485245",
		16#6057# => X"4144202d",
		16#6058# => X"444d554c",
		16#6059# => X"54495448",
		16#605a# => X"52454144",
		16#605b# => X"3d38202d",
		16#605c# => X"44504552",
		16#605d# => X"464f524d",
		16#605e# => X"414e4345",
		16#605f# => X"5f52554e",
		16#6060# => X"3d312020",
		16#6061# => X"2d6d6e65",
		16#6062# => X"776c6962",
		16#6063# => X"202d6d62",
		16#6064# => X"6f617264",
		16#6065# => X"3d6d6c35",
		16#6066# => X"30395f32",
		16#6067# => X"35005061",
		16#6068# => X"72616c6c",
		16#6069# => X"656c2025",
		16#606a# => X"73203a20",
		16#606b# => X"25640a00",
		16#606c# => X"50617261",
		16#606d# => X"4e757420",
		16#606e# => X"54687265",
		16#606f# => X"61647300",
		16#6070# => X"4d656d6f",
		16#6071# => X"7279206c",
		16#6072# => X"6f636174",
		16#6073# => X"696f6e20",
		16#6074# => X"203a2025",
		16#6075# => X"730a0053",
		16#6076# => X"5441434b",
		16#6077# => X"00736565",
		16#6078# => X"64637263",
		16#6079# => X"20202020",
		16#607a# => X"20202020",
		16#607b# => X"20203a20",
		16#607c# => X"30782530",
		16#607d# => X"34780a00",
		16#607e# => X"5b25645d",
		16#607f# => X"6372636c",
		16#6080# => X"69737420",
		16#6081# => X"20202020",
		16#6082# => X"20203a20",
		16#6083# => X"30782530",
		16#6084# => X"34780a00",
		16#6085# => X"5b25645d",
		16#6086# => X"6372636d",
		16#6087# => X"61747269",
		16#6088# => X"78202020",
		16#6089# => X"20203a20",
		16#608a# => X"30782530",
		16#608b# => X"34780a00",
		16#608c# => X"5b25645d",
		16#608d# => X"63726373",
		16#608e# => X"74617465",
		16#608f# => X"20202020",
		16#6090# => X"20203a20",
		16#6091# => X"30782530",
		16#6092# => X"34780a00",
		16#6093# => X"5b25645d",
		16#6094# => X"63726366",
		16#6095# => X"696e616c",
		16#6096# => X"20202020",
		16#6097# => X"20203a20",
		16#6098# => X"30782530",
		16#6099# => X"34780a00",
		16#609a# => X"436f7272",
		16#609b# => X"65637420",
		16#609c# => X"6f706572",
		16#609d# => X"6174696f",
		16#609e# => X"6e207661",
		16#609f# => X"6c696461",
		16#60a0# => X"7465642e",
		16#60a1# => X"20536565",
		16#60a2# => X"20726561",
		16#60a3# => X"646d652e",
		16#60a4# => X"74787420",
		16#60a5# => X"666f7220",
		16#60a6# => X"72756e20",
		16#60a7# => X"616e6420",
		16#60a8# => X"7265706f",
		16#60a9# => X"7274696e",
		16#60aa# => X"67207275",
		16#60ab# => X"6c65732e",
		16#60ac# => X"00436f72",
		16#60ad# => X"654d6172",
		16#60ae# => X"6b20312e",
		16#60af# => X"30203a20",
		16#60b0# => X"2566202f",
		16#60b1# => X"20257320",
		16#60b2# => X"25730020",
		16#60b3# => X"2f202573",
		16#60b4# => X"00202f20",
		16#60b5# => X"25643a25",
		16#60b6# => X"73004572",
		16#60b7# => X"726f7273",
		16#60b8# => X"20646574",
		16#60b9# => X"65637465",
		16#60ba# => X"64004361",
		16#60bb# => X"6e6e6f74",
		16#60bc# => X"2076616c",
		16#60bd# => X"69646174",
		16#60be# => X"65206f70",
		16#60bf# => X"65726174",
		16#60c0# => X"696f6e20",
		16#60c1# => X"666f7220",
		16#60c2# => X"74686573",
		16#60c3# => X"65207365",
		16#60c4# => X"65642076",
		16#60c5# => X"616c7565",
		16#60c6# => X"732c2070",
		16#60c7# => X"6c656173",
		16#60c8# => X"6520636f",
		16#60c9# => X"6d706172",
		16#60ca# => X"65207769",
		16#60cb# => X"74682072",
		16#60cc# => X"6573756c",
		16#60cd# => X"7473206f",
		16#60ce# => X"6e206120",
		16#60cf# => X"6b6e6f77",
		16#60d0# => X"6e20706c",
		16#60d1# => X"6174666f",
		16#60d2# => X"726d2e00",
		16#60d3# => X"53746174",
		16#60d4# => X"69630048",
		16#60d5# => X"65617000",
		16#60d6# => X"53746163",
		16#60d7# => X"6b000000",
		16#60d8# => X"3ff00000",
		16#60d9# => X"00000000",
		16#60da# => X"00000000",
		16#60db# => X"00000000",
		16#60dc# => X"40240000",
		16#60dd# => X"00000000",
		16#60de# => X"d4b03340",
		16#60df# => X"6a79e714",
		16#60e0# => X"e3c10000",
		16#60e1# => X"be521199",
		16#60e2# => X"56081fd7",
		16#60e3# => X"07470000",
		16#60e4# => X"5e4739bf",
		16#60e5# => X"e5a48e3a",
		16#60e6# => X"8d840000",
		16#60e7# => X"00005aa4",
		16#60e8# => X"00005aa4",
		16#60e9# => X"00005ac4",
		16#60ea# => X"00005ac4",
		16#60eb# => X"00005ae4",
		16#60ec# => X"00005cc8",
		16#60ed# => X"00005cb8",
		16#60ee# => X"00005c58",
		16#60ef# => X"00005d10",
		16#60f0# => X"00005c84",
		16#60f1# => X"00005c0c",
		16#60f2# => X"00005bb0",
		16#60f3# => X"00005b74",
		16#60f4# => X"00018410",
		16#60f5# => X"00018415",
		16#60f6# => X"0001841a",
		16#60f7# => X"0001841f",
		16#60f8# => X"00018424",
		16#60f9# => X"0001842d",
		16#60fa# => X"00018436",
		16#60fb# => X"0001843f",
		16#60fc# => X"00018448",
		16#60fd# => X"00018451",
		16#60fe# => X"0001845a",
		16#60ff# => X"00018463",
		16#6100# => X"0001846c",
		16#6101# => X"00018475",
		16#6102# => X"0001847e",
		16#6103# => X"00018487",
		16#6104# => X"35303132",
		16#6105# => X"00313233",
		16#6106# => X"34002d38",
		16#6107# => X"3734002b",
		16#6108# => X"31323200",
		16#6109# => X"33352e35",
		16#610a# => X"34343030",
		16#610b# => X"002e3132",
		16#610c# => X"33343530",
		16#610d# => X"30002d31",
		16#610e# => X"31302e37",
		16#610f# => X"3030002b",
		16#6110# => X"302e3634",
		16#6111# => X"34303000",
		16#6112# => X"352e3530",
		16#6113# => X"30652b33",
		16#6114# => X"002d2e31",
		16#6115# => X"3233652d",
		16#6116# => X"32002d38",
		16#6117# => X"37652b38",
		16#6118# => X"3332002b",
		16#6119# => X"302e3665",
		16#611a# => X"2d313200",
		16#611b# => X"54302e33",
		16#611c# => X"652d3146",
		16#611d# => X"002d542e",
		16#611e# => X"542b2b54",
		16#611f# => X"71003154",
		16#6120# => X"332e3465",
		16#6121# => X"347a0033",
		16#6122# => X"342e3065",
		16#6123# => X"2d545e00",
		16#6124# => X"000060dc",
		16#6125# => X"00006108",
		16#6126# => X"00006120",
		16#6127# => X"00006138",
		16#6128# => X"00006150",
		16#6129# => X"00006168",
		16#612a# => X"4572726f",
		16#612b# => X"7220616c",
		16#612c# => X"6c6f6361",
		16#612d# => X"74696e67",
		16#612e# => X"206d656d",
		16#612f# => X"6f727900",
		16#6130# => X"52756e6e",
		16#6131# => X"696e6720",
		16#6132# => X"436f7265",
		16#6133# => X"4d61726b",
		16#6134# => X"20776974",
		16#6135# => X"68202564",
		16#6136# => X"20636f72",
		16#6137# => X"65287329",
		16#6138# => X"2e2e2e0a",
		16#6139# => X"00000000",
		16#613a# => X"408f4000",
		16#613b# => X"00000000",
		16#613c# => X"28637075",
		16#613d# => X"69642023",
		16#613e# => X"25642920",
		16#613f# => X"2d2d2d2d",
		16#6140# => X"2d2d2d2d",
		16#6141# => X"2d2d2d2d",
		16#6142# => X"2d2d2d2d",
		16#6143# => X"2d2d2d2d",
		16#6144# => X"2d2d2d2d",
		16#6145# => X"2d2d2d2d",
		16#6146# => X"2d2d2d2d",
		16#6147# => X"2d2d2d2d",
		16#6148# => X"2d2d2d2d",
		16#6149# => X"2d2d2d2d",
		16#614a# => X"2d2d2d2d",
		16#614b# => X"2d2d2d2d",
		16#614c# => X"2d2d2d2d",
		16#614d# => X"2d2d2d2d",
		16#614e# => X"2d2d0a00",
		16#614f# => X"28637075",
		16#6150# => X"69642023",
		16#6151# => X"25642920",
		16#6152# => X"50657266",
		16#6153# => X"6f726d61",
		16#6154# => X"6e636520",
		16#6155# => X"73746174",
		16#6156# => X"69737469",
		16#6157# => X"63730a00",
		16#6158# => X"28637075",
		16#6159# => X"69642023",
		16#615a# => X"25642920",
		16#615b# => X"25377325",
		16#615c# => X"31317325",
		16#615d# => X"34732538",
		16#615e# => X"73253873",
		16#615f# => X"25313273",
		16#6160# => X"25313073",
		16#6161# => X"0a004576",
		16#6162# => X"656e7400",
		16#6163# => X"436f756e",
		16#6164# => X"74006d69",
		16#6165# => X"6e006176",
		16#6166# => X"67006d61",
		16#6167# => X"7800546f",
		16#6168# => X"74616c00",
		16#6169# => X"52617465",
		16#616a# => X"00286370",
		16#616b# => X"75696420",
		16#616c# => X"23256429",
		16#616d# => X"20253773",
		16#616e# => X"25313175",
		16#616f# => X"25347525",
		16#6170# => X"382e3266",
		16#6171# => X"25387525",
		16#6172# => X"31327525",
		16#6173# => X"31302e35",
		16#6174# => X"660a0041",
		16#6175# => X"4c550053",
		16#6176# => X"48494654",
		16#6177# => X"004d554c",
		16#6178# => X"004a554d",
		16#6179# => X"50004f54",
		16#617a# => X"48455200",
		16#617b# => X"28637075",
		16#617c# => X"69642023",
		16#617d# => X"25642920",
		16#617e# => X"25377325",
		16#617f# => X"31317525",
		16#6180# => X"34752538",
		16#6181# => X"2e326625",
		16#6182# => X"38752531",
		16#6183# => X"32750a00",
		16#6184# => X"414c4c00",
		16#6185# => X"43524849",
		16#6186# => X"46550043",
		16#6187# => X"524d4946",
		16#6188# => X"55004352",
		16#6189# => X"484c5355",
		16#618a# => X"0043524d",
		16#618b# => X"4c535500",
		16#618c# => X"4357484c",
		16#618d# => X"53550043",
		16#618e# => X"574d4c53",
		16#618f# => X"55002820",
		16#6190# => X"676c6f62",
		16#6191# => X"616c2029",
		16#6192# => X"202d2d2d",
		16#6193# => X"2d2d2d2d",
		16#6194# => X"2d2d2d2d",
		16#6195# => X"2d2d2d2d",
		16#6196# => X"2d2d2d2d",
		16#6197# => X"2d2d2d2d",
		16#6198# => X"2d2d2d2d",
		16#6199# => X"2d2d2d2d",
		16#619a# => X"2d2d2d2d",
		16#619b# => X"2d2d2d2d",
		16#619c# => X"2d2d2d2d",
		16#619d# => X"2d2d2d2d",
		16#619e# => X"2d2d2d2d",
		16#619f# => X"2d2d2d2d",
		16#61a0# => X"2d2d2d2d",
		16#61a1# => X"2d2d2d00",
		16#61a2# => X"2820676c",
		16#61a3# => X"6f62616c",
		16#61a4# => X"20292047",
		16#61a5# => X"6c6f6261",
		16#61a6# => X"6c207065",
		16#61a7# => X"72666f72",
		16#61a8# => X"6d616e63",
		16#61a9# => X"65207374",
		16#61aa# => X"61746973",
		16#61ab# => X"74696373",
		16#61ac# => X"00282067",
		16#61ad# => X"6c6f6261",
		16#61ae# => X"6c202920",
		16#61af# => X"25377325",
		16#61b0# => X"31317325",
		16#61b1# => X"34732538",
		16#61b2# => X"73253873",
		16#61b3# => X"25313273",
		16#61b4# => X"25313073",
		16#61b5# => X"0a002820",
		16#61b6# => X"676c6f62",
		16#61b7# => X"616c2029",
		16#61b8# => X"20253773",
		16#61b9# => X"25313175",
		16#61ba# => X"25347525",
		16#61bb# => X"382e3266",
		16#61bc# => X"25387525",
		16#61bd# => X"31327525",
		16#61be# => X"31302e35",
		16#61bf# => X"660a0028",
		16#61c0# => X"20676c6f",
		16#61c1# => X"62616c20",
		16#61c2# => X"29202537",
		16#61c3# => X"73253131",
		16#61c4# => X"75253475",
		16#61c5# => X"25382e32",
		16#61c6# => X"66253875",
		16#61c7# => X"25313275",
		16#61c8# => X"0a00434c",
		16#61c9# => X"4600434c",
		16#61ca# => X"57420028",
		16#61cb# => X"63707569",
		16#61cc# => X"64202325",
		16#61cd# => X"64292025",
		16#61ce# => X"735b2532",
		16#61cf# => X"645d2020",
		16#61d0# => X"20202020",
		16#61d1# => X"3a202564",
		16#61d2# => X"0a00696e",
		16#61d3# => X"736e204c",
		16#61d4# => X"4f414400",
		16#61d5# => X"696e736e",
		16#61d6# => X"2053544f",
		16#61d7# => X"52450000",
		16#61d8# => X"41e00000",
		16#61d9# => X"00000000",
		16#61da# => X"cf000000",
		16#61db# => X"00000000",
		16#61dc# => X"00000000",
		16#61dd# => X"00000000",
		16#61de# => X"00000000",
		16#61df# => X"00000000",
		16#61e0# => X"00000000",
		16#61e1# => X"00000000",
		16#61e2# => X"00000000",
		16#61e3# => X"00000000",
		16#61e4# => X"00010202",
		16#61e5# => X"03030303",
		16#61e6# => X"04040404",
		16#61e7# => X"04040404",
		16#61e8# => X"05050505",
		16#61e9# => X"05050505",
		16#61ea# => X"05050505",
		16#61eb# => X"05050505",
		16#61ec# => X"06060606",
		16#61ed# => X"06060606",
		16#61ee# => X"06060606",
		16#61ef# => X"06060606",
		16#61f0# => X"06060606",
		16#61f1# => X"06060606",
		16#61f2# => X"06060606",
		16#61f3# => X"06060606",
		16#61f4# => X"07070707",
		16#61f5# => X"07070707",
		16#61f6# => X"07070707",
		16#61f7# => X"07070707",
		16#61f8# => X"07070707",
		16#61f9# => X"07070707",
		16#61fa# => X"07070707",
		16#61fb# => X"07070707",
		16#61fc# => X"07070707",
		16#61fd# => X"07070707",
		16#61fe# => X"07070707",
		16#61ff# => X"07070707",
		16#6200# => X"07070707",
		16#6201# => X"07070707",
		16#6202# => X"07070707",
		16#6203# => X"07070707",
		16#6204# => X"08080808",
		16#6205# => X"08080808",
		16#6206# => X"08080808",
		16#6207# => X"08080808",
		16#6208# => X"08080808",
		16#6209# => X"08080808",
		16#620a# => X"08080808",
		16#620b# => X"08080808",
		16#620c# => X"08080808",
		16#620d# => X"08080808",
		16#620e# => X"08080808",
		16#620f# => X"08080808",
		16#6210# => X"08080808",
		16#6211# => X"08080808",
		16#6212# => X"08080808",
		16#6213# => X"08080808",
		16#6214# => X"08080808",
		16#6215# => X"08080808",
		16#6216# => X"08080808",
		16#6217# => X"08080808",
		16#6218# => X"08080808",
		16#6219# => X"08080808",
		16#621a# => X"08080808",
		16#621b# => X"08080808",
		16#621c# => X"08080808",
		16#621d# => X"08080808",
		16#621e# => X"08080808",
		16#621f# => X"08080808",
		16#6220# => X"08080808",
		16#6221# => X"08080808",
		16#6222# => X"08080808",
		16#6223# => X"08080808",
		16#6224# => X"0001ade8",
		16#6225# => X"4300494e",
		16#6226# => X"4600696e",
		16#6227# => X"66004e41",
		16#6228# => X"4e006e61",
		16#6229# => X"6e003031",
		16#622a# => X"32333435",
		16#622b# => X"36373839",
		16#622c# => X"41424344",
		16#622d# => X"45460030",
		16#622e# => X"31323334",
		16#622f# => X"35363738",
		16#6230# => X"39616263",
		16#6231# => X"64656600",
		16#6232# => X"286e756c",
		16#6233# => X"6c290000",
		16#6234# => X"00000000",
		16#6235# => X"00000000",
		16#6236# => X"0000e2d4",
		16#6237# => X"0000dd48",
		16#6238# => X"0000dd48",
		16#6239# => X"0000e2e8",
		16#623a# => X"0000dd48",
		16#623b# => X"0000dd48",
		16#623c# => X"0000dd48",
		16#623d# => X"0000dd48",
		16#623e# => X"0000dd48",
		16#623f# => X"0000dd48",
		16#6240# => X"0000deb0",
		16#6241# => X"0000e2f8",
		16#6242# => X"0000dd48",
		16#6243# => X"0000ded8",
		16#6244# => X"0000e344",
		16#6245# => X"0000dd48",
		16#6246# => X"0000e300",
		16#6247# => X"0000e310",
		16#6248# => X"0000e310",
		16#6249# => X"0000e310",
		16#624a# => X"0000e310",
		16#624b# => X"0000e310",
		16#624c# => X"0000e310",
		16#624d# => X"0000e310",
		16#624e# => X"0000e310",
		16#624f# => X"0000e310",
		16#6250# => X"0000dd48",
		16#6251# => X"0000dd48",
		16#6252# => X"0000dd48",
		16#6253# => X"0000dd48",
		16#6254# => X"0000dd48",
		16#6255# => X"0000dd48",
		16#6256# => X"0000dd48",
		16#6257# => X"0000dd48",
		16#6258# => X"0000dd48",
		16#6259# => X"0000dd48",
		16#625a# => X"0000e054",
		16#625b# => X"0000e180",
		16#625c# => X"0000dd48",
		16#625d# => X"0000e180",
		16#625e# => X"0000dd48",
		16#625f# => X"0000dd48",
		16#6260# => X"0000dd48",
		16#6261# => X"0000dd48",
		16#6262# => X"0000e260",
		16#6263# => X"0000dd48",
		16#6264# => X"0000dd48",
		16#6265# => X"0000e5fc",
		16#6266# => X"0000dd48",
		16#6267# => X"0000dd48",
		16#6268# => X"0000dd48",
		16#6269# => X"0000dd48",
		16#626a# => X"0000dd48",
		16#626b# => X"0000e564",
		16#626c# => X"0000dd48",
		16#626d# => X"0000dd48",
		16#626e# => X"0000e5ac",
		16#626f# => X"0000dd48",
		16#6270# => X"0000dd48",
		16#6271# => X"0000dd48",
		16#6272# => X"0000dd48",
		16#6273# => X"0000dd48",
		16#6274# => X"0000dd48",
		16#6275# => X"0000dd48",
		16#6276# => X"0000dd48",
		16#6277# => X"0000dd48",
		16#6278# => X"0000dd48",
		16#6279# => X"0000e270",
		16#627a# => X"0000e2a8",
		16#627b# => X"0000e180",
		16#627c# => X"0000e180",
		16#627d# => X"0000e180",
		16#627e# => X"0000e39c",
		16#627f# => X"0000e2a8",
		16#6280# => X"0000dd48",
		16#6281# => X"0000dd48",
		16#6282# => X"0000e3ac",
		16#6283# => X"0000dd48",
		16#6284# => X"0000e3bc",
		16#6285# => X"0000e644",
		16#6286# => X"0000e3f0",
		16#6287# => X"0000e554",
		16#6288# => X"0000dd48",
		16#6289# => X"0000e450",
		16#628a# => X"0000dd48",
		16#628b# => X"0000e64c",
		16#628c# => X"0000dd48",
		16#628d# => X"0000dd48",
		16#628e# => X"0000e4c4",
		16#628f# => X"30303030",
		16#6290# => X"30303030",
		16#6291# => X"30303030",
		16#6292# => X"30303030",
		16#6293# => X"20202020",
		16#6294# => X"20202020",
		16#6295# => X"20202020",
		16#6296# => X"20202020",
		16#6297# => X"496e6669",
		16#6298# => X"6e697479",
		16#6299# => X"004e614e",
		16#629a# => X"00000000",
		16#629b# => X"00000000",
		16#629c# => X"00000000",
		16#629d# => X"3ff80000",
		16#629e# => X"00000000",
		16#629f# => X"3fd287a7",
		16#62a0# => X"636f4361",
		16#62a1# => X"3fc68a28",
		16#62a2# => X"8b60c8b3",
		16#62a3# => X"3fd34413",
		16#62a4# => X"509f79fb",
		16#62a5# => X"3ff00000",
		16#62a6# => X"00000000",
		16#62a7# => X"40240000",
		16#62a8# => X"00000000",
		16#62a9# => X"401c0000",
		16#62aa# => X"00000000",
		16#62ab# => X"40140000",
		16#62ac# => X"00000000",
		16#62ad# => X"3fe00000",
		16#62ae# => X"00000000",
		16#62af# => X"504f5349",
		16#62b0# => X"58000000",
		16#62b1# => X"00017f76",
		16#62b2# => X"0001853b",
		16#62b3# => X"0001853b",
		16#62b4# => X"0001853b",
		16#62b5# => X"0001853b",
		16#62b6# => X"0001853b",
		16#62b7# => X"0001853b",
		16#62b8# => X"0001853b",
		16#62b9# => X"0001853b",
		16#62ba# => X"0001853b",
		16#62bb# => X"7f7f7f7f",
		16#62bc# => X"7f7f7f7f",
		16#62bd# => X"7f7f7f7f",
		16#62be# => X"7f7f0000",
		16#62bf# => X"40240000",
		16#62c0# => X"00000000",
		16#62c1# => X"3ff00000",
		16#62c2# => X"00000000",
		16#62c3# => X"40240000",
		16#62c4# => X"00000000",
		16#62c5# => X"40590000",
		16#62c6# => X"00000000",
		16#62c7# => X"408f4000",
		16#62c8# => X"00000000",
		16#62c9# => X"40c38800",
		16#62ca# => X"00000000",
		16#62cb# => X"40f86a00",
		16#62cc# => X"00000000",
		16#62cd# => X"412e8480",
		16#62ce# => X"00000000",
		16#62cf# => X"416312d0",
		16#62d0# => X"00000000",
		16#62d1# => X"4197d784",
		16#62d2# => X"00000000",
		16#62d3# => X"41cdcd65",
		16#62d4# => X"00000000",
		16#62d5# => X"4202a05f",
		16#62d6# => X"20000000",
		16#62d7# => X"42374876",
		16#62d8# => X"e8000000",
		16#62d9# => X"426d1a94",
		16#62da# => X"a2000000",
		16#62db# => X"42a2309c",
		16#62dc# => X"e5400000",
		16#62dd# => X"42d6bcc4",
		16#62de# => X"1e900000",
		16#62df# => X"430c6bf5",
		16#62e0# => X"26340000",
		16#62e1# => X"4341c379",
		16#62e2# => X"37e08000",
		16#62e3# => X"43763457",
		16#62e4# => X"85d8a000",
		16#62e5# => X"43abc16d",
		16#62e6# => X"674ec800",
		16#62e7# => X"43e158e4",
		16#62e8# => X"60913d00",
		16#62e9# => X"4415af1d",
		16#62ea# => X"78b58c40",
		16#62eb# => X"444b1ae4",
		16#62ec# => X"d6e2ef50",
		16#62ed# => X"4480f0cf",
		16#62ee# => X"064dd592",
		16#62ef# => X"44b52d02",
		16#62f0# => X"c7e14af6",
		16#62f1# => X"44ea7843",
		16#62f2# => X"79d99db4",
		16#62f3# => X"4341c379",
		16#62f4# => X"37e08000",
		16#62f5# => X"4693b8b5",
		16#62f6# => X"b5056e17",
		16#62f7# => X"4d384f03",
		16#62f8# => X"e93ff9f5",
		16#62f9# => X"5a827748",
		16#62fa# => X"f9301d32",
		16#62fb# => X"75154fdd",
		16#62fc# => X"7f73bf3c",
		16#62fd# => X"3c9cd2b2",
		16#62fe# => X"97d889bc",
		16#62ff# => X"3949f623",
		16#6300# => X"d5a8a733",
		16#6301# => X"32a50ffd",
		16#6302# => X"44f4a73d",
		16#6303# => X"255bba08",
		16#6304# => X"cf8c979d",
		16#6305# => X"0ac80628",
		16#6306# => X"64ac6f43",
		16#6307# => X"00000005",
		16#6308# => X"00000019",
		16#6309# => X"0000007d",
		16#630a# => X"000163e4",
		16#630b# => X"00015f54",
		16#630c# => X"00015f54",
		16#630d# => X"000163dc",
		16#630e# => X"00015f54",
		16#630f# => X"00015f54",
		16#6310# => X"00015f54",
		16#6311# => X"00015f54",
		16#6312# => X"00015f54",
		16#6313# => X"00015f54",
		16#6314# => X"000161d8",
		16#6315# => X"00016208",
		16#6316# => X"00015f54",
		16#6317# => X"00016200",
		16#6318# => X"00016218",
		16#6319# => X"00015f54",
		16#631a# => X"00016210",
		16#631b# => X"000164a0",
		16#631c# => X"000164a0",
		16#631d# => X"000164a0",
		16#631e# => X"000164a0",
		16#631f# => X"000164a0",
		16#6320# => X"000164a0",
		16#6321# => X"000164a0",
		16#6322# => X"000164a0",
		16#6323# => X"000164a0",
		16#6324# => X"00015f54",
		16#6325# => X"00015f54",
		16#6326# => X"00015f54",
		16#6327# => X"00015f54",
		16#6328# => X"00015f54",
		16#6329# => X"00015f54",
		16#632a# => X"00015f54",
		16#632b# => X"00015f54",
		16#632c# => X"00015f54",
		16#632d# => X"00015f54",
		16#632e# => X"00016494",
		16#632f# => X"00015f54",
		16#6330# => X"00015f54",
		16#6331# => X"00015f54",
		16#6332# => X"00015f54",
		16#6333# => X"00015f54",
		16#6334# => X"00015f54",
		16#6335# => X"00015f54",
		16#6336# => X"00015f54",
		16#6337# => X"00015f54",
		16#6338# => X"00015f54",
		16#6339# => X"000160a0",
		16#633a# => X"00015f54",
		16#633b# => X"00015f54",
		16#633c# => X"00015f54",
		16#633d# => X"00015f54",
		16#633e# => X"00015f54",
		16#633f# => X"0001619c",
		16#6340# => X"00015f54",
		16#6341# => X"00015f54",
		16#6342# => X"00016480",
		16#6343# => X"00015f54",
		16#6344# => X"00015f54",
		16#6345# => X"00015f54",
		16#6346# => X"00015f54",
		16#6347# => X"00015f54",
		16#6348# => X"00015f54",
		16#6349# => X"00015f54",
		16#634a# => X"00015f54",
		16#634b# => X"00015f54",
		16#634c# => X"00015f54",
		16#634d# => X"00016450",
		16#634e# => X"00016400",
		16#634f# => X"00015f54",
		16#6350# => X"00015f54",
		16#6351# => X"00015f54",
		16#6352# => X"000163f8",
		16#6353# => X"00016400",
		16#6354# => X"00015f54",
		16#6355# => X"00015f54",
		16#6356# => X"00016098",
		16#6357# => X"00015f54",
		16#6358# => X"00016270",
		16#6359# => X"000160a4",
		16#635a# => X"00016330",
		16#635b# => X"00016098",
		16#635c# => X"00015f54",
		16#635d# => X"00016378",
		16#635e# => X"00015f54",
		16#635f# => X"000161a0",
		16#6360# => X"00015f54",
		16#6361# => X"00015f54",
		16#6362# => X"000162a8",
		16#6363# => X"30303030",
		16#6364# => X"30303030",
		16#6365# => X"30303030",
		16#6366# => X"30303030",
		16#6367# => X"20202020",
		16#6368# => X"20202020",
		16#6369# => X"20202020",
		16#636a# => X"20202020",
		16#636b# => X"00000000",
		16#636c# => X"00000000",
		16#636d# => X"00000000",
		16#636e# => X"00000000",
		16#636f# => X"00000000",
		16#6370# => X"00000000",
		16#6371# => X"00000000",
		16#6372# => X"00000000",
		16#6373# => X"00000000",
		16#6374# => X"00000000",
		16#6375# => X"00000000",
		16#6376# => X"00000000",
		16#6377# => X"00000000",
		16#6378# => X"00000000",
		16#6379# => X"00000000",
		16#637a# => X"00000000",
		16#637b# => X"00000000",
		16#637c# => X"00000000",
		16#637d# => X"00000000",
		16#637e# => X"00000000",
		16#637f# => X"00000000",
		16#6380# => X"00000000",
		16#6381# => X"00000000",
		16#6382# => X"00000000",
		16#6383# => X"00000000",
		16#6384# => X"00000000",
		16#6385# => X"00000000",
		16#6386# => X"00000000",
		16#6387# => X"00000000",
		16#6388# => X"00000000",
		16#6389# => X"00000000",
		16#638a# => X"00000000",
		16#638b# => X"00000000",
		16#638c# => X"00000000",
		16#638d# => X"00000000",
		16#638e# => X"00000000",
		16#638f# => X"00000000",
		16#6390# => X"00000000",
		16#6391# => X"00000000",
		16#6392# => X"00000000",
		16#6393# => X"00000000",
		16#6394# => X"00000000",
		16#6395# => X"00000000",
		16#6396# => X"00000000",
		16#6397# => X"00000000",
		16#6398# => X"00000000",
		16#6399# => X"00000000",
		16#639a# => X"00000000",
		16#639b# => X"00000000",
		16#639c# => X"00000000",
		16#639d# => X"00000000",
		16#639e# => X"00000000",
		16#639f# => X"00000000",
		16#63a0# => X"00000000",
		16#63a1# => X"00000000",
		16#63a2# => X"00000000",
		16#63a3# => X"00000000",
		16#63a4# => X"00000000",
		16#63a5# => X"00000000",
		16#63a6# => X"00000000",
		16#63a7# => X"00000000",
		16#63a8# => X"00000000",
		16#63a9# => X"00000000",
		16#63aa# => X"00000000",
		16#63ab# => X"00000000",
		16#63ac# => X"00000000",
		16#63ad# => X"00000000",
		16#63ae# => X"00000000",
		16#63af# => X"00000000",
		16#63b0# => X"00000000",
		16#63b1# => X"00000000",
		16#63b2# => X"00000000",
		16#63b3# => X"00000000",
		16#63b4# => X"00000000",
		16#63b5# => X"00000000",
		16#63b6# => X"00000000",
		16#63b7# => X"00000000",
		16#63b8# => X"00000000",
		16#63b9# => X"00000000",
		16#63ba# => X"00000000",
		16#63bb# => X"00000000",
		16#63bc# => X"00000000",
		16#63bd# => X"00000000",
		16#63be# => X"00000000",
		16#63bf# => X"00000000",
		16#63c0# => X"00000000",
		16#63c1# => X"00000000",
		16#63c2# => X"00000000",
		16#63c3# => X"00000000",
		16#63c4# => X"00000000",
		16#63c5# => X"00000000",
		16#63c6# => X"00000000",
		16#63c7# => X"00000000",
		16#63c8# => X"00000000",
		16#63c9# => X"00000000",
		16#63ca# => X"00000000",
		16#63cb# => X"00000000",
		16#63cc# => X"00000000",
		16#63cd# => X"00000000",
		16#63ce# => X"00000000",
		16#63cf# => X"00000000",
		16#63d0# => X"00000000",
		16#63d1# => X"00000000",
		16#63d2# => X"00000000",
		16#63d3# => X"00000000",
		16#63d4# => X"00000000",
		16#63d5# => X"00000000",
		16#63d6# => X"00000000",
		16#63d7# => X"00000000",
		16#63d8# => X"00000000",
		16#63d9# => X"00000000",
		16#63da# => X"00000000",
		16#63db# => X"00000000",
		16#63dc# => X"00000000",
		16#63dd# => X"00000000",
		16#63de# => X"00000000",
		16#63df# => X"00000000",
		16#63e0# => X"00000000",
		16#63e1# => X"00000000",
		16#63e2# => X"00000000",
		16#63e3# => X"00000000",
		16#63e4# => X"00000000",
		16#63e5# => X"00000000",
		16#63e6# => X"00000000",
		16#63e7# => X"00000000",
		16#63e8# => X"00000000",
		16#63e9# => X"00000000",
		16#63ea# => X"00000000",
		16#63eb# => X"00000000",
		16#63ec# => X"00000000",
		16#63ed# => X"00000000",
		16#63ee# => X"00000000",
		16#63ef# => X"00000000",
		16#63f0# => X"00000000",
		16#63f1# => X"00000000",
		16#63f2# => X"00000000",
		16#63f3# => X"00000000",
		16#63f4# => X"00000000",
		16#63f5# => X"00000000",
		16#63f6# => X"00000000",
		16#63f7# => X"00000000",
		16#63f8# => X"00000000",
		16#63f9# => X"00000000",
		16#63fa# => X"00000000",
		16#63fb# => X"00000000",
		16#63fc# => X"00000000",
		16#63fd# => X"00000000",
		16#63fe# => X"00000000",
		16#63ff# => X"00000000",
		16#6400# => X"00000000",
		16#6401# => X"00000000",
		16#6402# => X"00000000",
		16#6403# => X"00000000",
		16#6404# => X"00000000",
		16#6405# => X"00000000",
		16#6406# => X"00000000",
		16#6407# => X"00000000",
		16#6408# => X"00000000",
		16#6409# => X"00000000",
		16#640a# => X"00000000",
		16#640b# => X"00000000",
		16#640c# => X"00000000",
		16#640d# => X"00000000",
		16#640e# => X"00000000",
		16#640f# => X"00000000",
		16#6410# => X"00000000",
		16#6411# => X"00000000",
		16#6412# => X"00000000",
		16#6413# => X"00000000",
		16#6414# => X"00000000",
		16#6415# => X"00000000",
		16#6416# => X"00000000",
		16#6417# => X"00000000",
		16#6418# => X"00000000",
		16#6419# => X"00000000",
		16#641a# => X"00000000",
		16#641b# => X"00000000",
		16#641c# => X"00000000",
		16#641d# => X"00000000",
		16#641e# => X"00000000",
		16#641f# => X"00000000",
		16#6420# => X"00000000",
		16#6421# => X"00000000",
		16#6422# => X"00000000",
		16#6423# => X"00000000",
		16#6424# => X"00000000",
		16#6425# => X"00000000",
		16#6426# => X"00000000",
		16#6427# => X"00000000",
		16#6428# => X"00000000",
		16#6429# => X"00000000",
		16#642a# => X"00000000",
		16#642b# => X"00000000",
		16#642c# => X"00000000",
		16#642d# => X"00000000",
		16#642e# => X"00000000",
		16#642f# => X"00000000",
		16#6430# => X"00000000",
		16#6431# => X"00000000",
		16#6432# => X"00000000",
		16#6433# => X"00000000",
		16#6434# => X"00000000",
		16#6435# => X"00000000",
		16#6436# => X"00000000",
		16#6437# => X"00000000",
		16#6438# => X"00000000",
		16#6439# => X"00000000",
		16#643a# => X"00000000",
		16#643b# => X"00000000",
		16#643c# => X"00000000",
		16#643d# => X"00000000",
		16#643e# => X"00000000",
		16#643f# => X"00000000",
		16#6440# => X"00000000",
		16#6441# => X"00000000",
		16#6442# => X"00000000",
		16#6443# => X"00000000",
		16#6444# => X"00000000",
		16#6445# => X"00000000",
		16#6446# => X"00000000",
		16#6447# => X"00000000",
		16#6448# => X"00000000",
		16#6449# => X"00000000",
		16#644a# => X"00000000",
		16#644b# => X"00000000",
		16#644c# => X"00000000",
		16#644d# => X"00000000",
		16#644e# => X"00000000",
		16#644f# => X"00000000",
		16#6450# => X"00000000",
		16#6451# => X"00000000",
		16#6452# => X"00000000",
		16#6453# => X"00000000",
		16#6454# => X"00000000",
		16#6455# => X"00000000",
		16#6456# => X"00000000",
		16#6457# => X"00000000",
		16#6458# => X"00000000",
		16#6459# => X"00000000",
		16#645a# => X"00000000",
		16#645b# => X"00000000",
		16#645c# => X"00000000",
		16#645d# => X"00000000",
		16#645e# => X"00000000",
		16#645f# => X"00000000",
		16#6460# => X"00000000",
		16#6461# => X"00000000",
		16#6462# => X"00000000",
		16#6463# => X"00000000",
		16#6464# => X"00000000",
		16#6465# => X"00000000",
		16#6466# => X"00000000",
		16#6467# => X"00000000",
		16#6468# => X"00000000",
		16#6469# => X"00000000",
		16#646a# => X"00000000",
		16#646b# => X"00000000",
		16#646c# => X"00000000",
		16#646d# => X"00000000",
		16#646e# => X"00000000",
		16#646f# => X"00000000",
		16#6470# => X"00000000",
		16#6471# => X"00000000",
		16#6472# => X"00000000",
		16#6473# => X"00000000",
		16#6474# => X"00000000",
		16#6475# => X"00000000",
		16#6476# => X"00000000",
		16#6477# => X"00000000",
		16#6478# => X"00000000",
		16#6479# => X"00000000",
		16#647a# => X"00000000",
		16#647b# => X"00000000",
		16#647c# => X"00000000",
		16#647d# => X"00000000",
		16#647e# => X"00000000",
		16#647f# => X"00000000",
		16#6480# => X"00000000",
		16#6481# => X"00000000",
		16#6482# => X"00000000",
		16#6483# => X"00000000",
		16#6484# => X"00000000",
		16#6485# => X"00000000",
		16#6486# => X"00000000",
		16#6487# => X"00000000",
		16#6488# => X"00000000",
		16#6489# => X"00000000",
		16#648a# => X"00000000",
		16#648b# => X"00000000",
		16#648c# => X"00000000",
		16#648d# => X"00000000",
		16#648e# => X"00000000",
		16#648f# => X"00000000",
		16#6490# => X"00000000",
		16#6491# => X"00000000",
		16#6492# => X"00000000",
		16#6493# => X"00000000",
		16#6494# => X"00000000",
		16#6495# => X"00000000",
		16#6496# => X"00000000",
		16#6497# => X"00000000",
		16#6498# => X"00000000",
		16#6499# => X"00000000",
		16#649a# => X"00000000",
		16#649b# => X"00000000",
		16#649c# => X"00000000",
		16#649d# => X"00000000",
		16#649e# => X"00000000",
		16#649f# => X"00000000",
		16#64a0# => X"00000000",
		16#64a1# => X"00000000",
		16#64a2# => X"00000000",
		16#64a3# => X"00000000",
		16#64a4# => X"00000000",
		16#64a5# => X"00000000",
		16#64a6# => X"00000000",
		16#64a7# => X"00000000",
		16#64a8# => X"00000000",
		16#64a9# => X"00000000",
		16#64aa# => X"00000000",
		16#64ab# => X"00000000",
		16#64ac# => X"00000000",
		16#64ad# => X"00000000",
		16#64ae# => X"00000000",
		16#64af# => X"00000000",
		16#64b0# => X"00000000",
		16#64b1# => X"00000000",
		16#64b2# => X"00000000",
		16#64b3# => X"00000000",
		16#64b4# => X"00000000",
		16#64b5# => X"00000000",
		16#64b6# => X"00000000",
		16#64b7# => X"00000000",
		16#64b8# => X"00000000",
		16#64b9# => X"00000000",
		16#64ba# => X"00000000",
		16#64bb# => X"00000000",
		16#64bc# => X"00000000",
		16#64bd# => X"00000000",
		16#64be# => X"00000000",
		16#64bf# => X"00000000",
		16#64c0# => X"00000000",
		16#64c1# => X"00000000",
		16#64c2# => X"00000000",
		16#64c3# => X"00000000",
		16#64c4# => X"00000000",
		16#64c5# => X"00000000",
		16#64c6# => X"00000000",
		16#64c7# => X"00000000",
		16#64c8# => X"00000000",
		16#64c9# => X"00000000",
		16#64ca# => X"00000000",
		16#64cb# => X"00000000",
		16#64cc# => X"00000000",
		16#64cd# => X"00000000",
		16#64ce# => X"00000000",
		16#64cf# => X"00000000",
		16#64d0# => X"00000000",
		16#64d1# => X"00000000",
		16#64d2# => X"00000000",
		16#64d3# => X"00000000",
		16#64d4# => X"00000000",
		16#64d5# => X"00000000",
		16#64d6# => X"00000000",
		16#64d7# => X"00000000",
		16#64d8# => X"00000000",
		16#64d9# => X"00000000",
		16#64da# => X"00000000",
		16#64db# => X"00000000",
		16#64dc# => X"00000000",
		16#64dd# => X"00000000",
		16#64de# => X"00000000",
		16#64df# => X"00000000",
		16#64e0# => X"00000000",
		16#64e1# => X"00000000",
		16#64e2# => X"00000000",
		16#64e3# => X"00000000",
		16#64e4# => X"00000000",
		16#64e5# => X"00000000",
		16#64e6# => X"00000000",
		16#64e7# => X"00000000",
		16#64e8# => X"00000000",
		16#64e9# => X"00000000",
		16#64ea# => X"00000000",
		16#64eb# => X"00000000",
		16#64ec# => X"00000000",
		16#64ed# => X"00000000",
		16#64ee# => X"00000000",
		16#64ef# => X"00000000",
		16#64f0# => X"00000000",
		16#64f1# => X"00000000",
		16#64f2# => X"00000000",
		16#64f3# => X"00000000",
		16#64f4# => X"00000000",
		16#64f5# => X"00000000",
		16#64f6# => X"00000000",
		16#64f7# => X"00000000",
		16#64f8# => X"00000000",
		16#64f9# => X"00000000",
		16#64fa# => X"00000000",
		16#64fb# => X"00000000",
		16#64fc# => X"00000000",
		16#64fd# => X"00000000",
		16#64fe# => X"00000000",
		16#64ff# => X"00000000",
		16#6500# => X"00000000",
		16#6501# => X"00000000",
		16#6502# => X"00000000",
		16#6503# => X"00000000",
		16#6504# => X"00000000",
		16#6505# => X"00000000",
		16#6506# => X"00000000",
		16#6507# => X"00000000",
		16#6508# => X"00000000",
		16#6509# => X"00000000",
		16#650a# => X"00000000",
		16#650b# => X"00000000",
		16#650c# => X"00000000",
		16#650d# => X"00000000",
		16#650e# => X"00000000",
		16#650f# => X"00000000",
		16#6510# => X"00000000",
		16#6511# => X"00000000",
		16#6512# => X"00000000",
		16#6513# => X"00000000",
		16#6514# => X"00000000",
		16#6515# => X"00000000",
		16#6516# => X"00000000",
		16#6517# => X"00000000",
		16#6518# => X"00000000",
		16#6519# => X"00000000",
		16#651a# => X"00000000",
		16#651b# => X"00000000",
		16#651c# => X"00000000",
		16#651d# => X"00000000",
		16#651e# => X"00000000",
		16#651f# => X"00000000",
		16#6520# => X"00000000",
		16#6521# => X"00000000",
		16#6522# => X"00000000",
		16#6523# => X"00000000",
		16#6524# => X"00000000",
		16#6525# => X"00000000",
		16#6526# => X"00000000",
		16#6527# => X"00000000",
		16#6528# => X"00000000",
		16#6529# => X"00000000",
		16#652a# => X"00000000",
		16#652b# => X"00000000",
		16#652c# => X"00000000",
		16#652d# => X"00000000",
		16#652e# => X"00000000",
		16#652f# => X"00000000",
		16#6530# => X"00000000",
		16#6531# => X"00000000",
		16#6532# => X"00000000",
		16#6533# => X"00000000",
		16#6534# => X"00000000",
		16#6535# => X"00000000",
		16#6536# => X"00000000",
		16#6537# => X"00000000",
		16#6538# => X"00000000",
		16#6539# => X"00000000",
		16#653a# => X"00000000",
		16#653b# => X"00000000",
		16#653c# => X"00000000",
		16#653d# => X"00000000",
		16#653e# => X"00000000",
		16#653f# => X"00000000",
		16#6540# => X"00000000",
		16#6541# => X"00000000",
		16#6542# => X"00000000",
		16#6543# => X"00000000",
		16#6544# => X"00000000",
		16#6545# => X"00000000",
		16#6546# => X"00000000",
		16#6547# => X"00000000",
		16#6548# => X"00000000",
		16#6549# => X"00000000",
		16#654a# => X"00000000",
		16#654b# => X"00000000",
		16#654c# => X"00000000",
		16#654d# => X"00000000",
		16#654e# => X"00000000",
		16#654f# => X"00000000",
		16#6550# => X"00000000",
		16#6551# => X"00000000",
		16#6552# => X"00000000",
		16#6553# => X"00000000",
		16#6554# => X"00000000",
		16#6555# => X"00000000",
		16#6556# => X"00000000",
		16#6557# => X"00000000",
		16#6558# => X"00000000",
		16#6559# => X"00000000",
		16#655a# => X"00000000",
		16#655b# => X"00000000",
		16#655c# => X"00000000",
		16#655d# => X"00000000",
		16#655e# => X"00000000",
		16#655f# => X"00000000",
		16#6560# => X"00000000",
		16#6561# => X"00000000",
		16#6562# => X"00000000",
		16#6563# => X"00000000",
		16#6564# => X"00000000",
		16#6565# => X"00000000",
		16#6566# => X"00000000",
		16#6567# => X"00000000",
		16#6568# => X"00000000",
		16#6569# => X"00000000",
		16#656a# => X"00000000",
		16#656b# => X"00000000",
		16#656c# => X"00000000",
		16#656d# => X"00000000",
		16#656e# => X"00000000",
		16#656f# => X"00000000",
		16#6570# => X"00000000",
		16#6571# => X"00000000",
		16#6572# => X"00000000",
		16#6573# => X"00000000",
		16#6574# => X"00000000",
		16#6575# => X"00000000",
		16#6576# => X"00000000",
		16#6577# => X"00000000",
		16#6578# => X"00000000",
		16#6579# => X"00000000",
		16#657a# => X"00000000",
		16#657b# => X"00000000",
		16#657c# => X"00000000",
		16#657d# => X"00000000",
		16#657e# => X"00000000",
		16#657f# => X"00000000",
		16#6580# => X"00000000",
		16#6581# => X"00000000",
		16#6582# => X"00000000",
		16#6583# => X"00000000",
		16#6584# => X"00000000",
		16#6585# => X"00000000",
		16#6586# => X"00000000",
		16#6587# => X"00000000",
		16#6588# => X"00000000",
		16#6589# => X"00000000",
		16#658a# => X"00000000",
		16#658b# => X"00000000",
		16#658c# => X"00000000",
		16#658d# => X"00000000",
		16#658e# => X"00000000",
		16#658f# => X"00000000",
		16#6590# => X"00000000",
		16#6591# => X"00000000",
		16#6592# => X"00000000",
		16#6593# => X"00000000",
		16#6594# => X"00000000",
		16#6595# => X"00000000",
		16#6596# => X"00000000",
		16#6597# => X"00000000",
		16#6598# => X"00000000",
		16#6599# => X"00000000",
		16#659a# => X"00000000",
		16#659b# => X"00000000",
		16#659c# => X"00000000",
		16#659d# => X"00000000",
		16#659e# => X"00000000",
		16#659f# => X"00000000",
		16#65a0# => X"00000000",
		16#65a1# => X"00000000",
		16#65a2# => X"00000000",
		16#65a3# => X"00000000",
		16#65a4# => X"00000000",
		16#65a5# => X"00000000",
		16#65a6# => X"00000000",
		16#65a7# => X"00000000",
		16#65a8# => X"00000000",
		16#65a9# => X"00000000",
		16#65aa# => X"00000000",
		16#65ab# => X"00000000",
		16#65ac# => X"00000000",
		16#65ad# => X"00000000",
		16#65ae# => X"00000000",
		16#65af# => X"00000000",
		16#65b0# => X"00000000",
		16#65b1# => X"00000000",
		16#65b2# => X"00000000",
		16#65b3# => X"00000000",
		16#65b4# => X"00000000",
		16#65b5# => X"00000000",
		16#65b6# => X"00000000",
		16#65b7# => X"00000000",
		16#65b8# => X"00000000",
		16#65b9# => X"00000000",
		16#65ba# => X"00000000",
		16#65bb# => X"00000000",
		16#65bc# => X"00000000",
		16#65bd# => X"00000000",
		16#65be# => X"00000000",
		16#65bf# => X"00000000",
		16#65c0# => X"00000000",
		16#65c1# => X"00000000",
		16#65c2# => X"00000000",
		16#65c3# => X"00000000",
		16#65c4# => X"00000000",
		16#65c5# => X"00000000",
		16#65c6# => X"00000000",
		16#65c7# => X"00000000",
		16#65c8# => X"00000000",
		16#65c9# => X"00000000",
		16#65ca# => X"00000000",
		16#65cb# => X"00000000",
		16#65cc# => X"00000000",
		16#65cd# => X"00000000",
		16#65ce# => X"00000000",
		16#65cf# => X"00000000",
		16#65d0# => X"00000000",
		16#65d1# => X"00000000",
		16#65d2# => X"00000000",
		16#65d3# => X"00000000",
		16#65d4# => X"00000000",
		16#65d5# => X"00000000",
		16#65d6# => X"00000000",
		16#65d7# => X"00000000",
		16#65d8# => X"00000000",
		16#65d9# => X"00000000",
		16#65da# => X"00000000",
		16#65db# => X"00000000",
		16#65dc# => X"00000000",
		16#65dd# => X"00000000",
		16#65de# => X"00000000",
		16#65df# => X"00000000",
		16#65e0# => X"00000000",
		16#65e1# => X"00000000",
		16#65e2# => X"00000000",
		16#65e3# => X"00000000",
		16#65e4# => X"00000000",
		16#65e5# => X"00000000",
		16#65e6# => X"00000000",
		16#65e7# => X"00000000",
		16#65e8# => X"00000000",
		16#65e9# => X"00000000",
		16#65ea# => X"00000000",
		16#65eb# => X"00000000",
		16#65ec# => X"00000000",
		16#65ed# => X"00000000",
		16#65ee# => X"00000000",
		16#65ef# => X"00000000",
		16#65f0# => X"00000000",
		16#65f1# => X"00000000",
		16#65f2# => X"00000000",
		16#65f3# => X"00000000",
		16#65f4# => X"00000000",
		16#65f5# => X"00000000",
		16#65f6# => X"00000000",
		16#65f7# => X"00000000",
		16#65f8# => X"00000000",
		16#65f9# => X"00000000",
		16#65fa# => X"00000000",
		16#65fb# => X"00000000",
		16#65fc# => X"00000000",
		16#65fd# => X"00000000",
		16#65fe# => X"00000000",
		16#65ff# => X"00000000",
		16#6600# => X"00000000",
		16#6601# => X"00000000",
		16#6602# => X"00000000",
		16#6603# => X"00000000",
		16#6604# => X"00000000",
		16#6605# => X"00000000",
		16#6606# => X"00000000",
		16#6607# => X"00000000",
		16#6608# => X"00000000",
		16#6609# => X"00000000",
		16#660a# => X"00000000",
		16#660b# => X"00000000",
		16#660c# => X"00000000",
		16#660d# => X"00000000",
		16#660e# => X"00000000",
		16#660f# => X"00000000",
		16#6610# => X"00000000",
		16#6611# => X"00000000",
		16#6612# => X"00000000",
		16#6613# => X"00000000",
		16#6614# => X"00000000",
		16#6615# => X"00000000",
		16#6616# => X"00000000",
		16#6617# => X"00000000",
		16#6618# => X"00000000",
		16#6619# => X"00000000",
		16#661a# => X"00000000",
		16#661b# => X"00000000",
		16#661c# => X"00000000",
		16#661d# => X"00000000",
		16#661e# => X"00000000",
		16#661f# => X"00000000",
		16#6620# => X"00000000",
		16#6621# => X"00000000",
		16#6622# => X"00000000",
		16#6623# => X"00000000",
		16#6624# => X"00000000",
		16#6625# => X"00000000",
		16#6626# => X"00000000",
		16#6627# => X"00000000",
		16#6628# => X"00000000",
		16#6629# => X"00000000",
		16#662a# => X"00000000",
		16#662b# => X"00000000",
		16#662c# => X"00000000",
		16#662d# => X"00000000",
		16#662e# => X"00000000",
		16#662f# => X"00000000",
		16#6630# => X"00000000",
		16#6631# => X"00000000",
		16#6632# => X"00000000",
		16#6633# => X"00000000",
		16#6634# => X"00000000",
		16#6635# => X"00000000",
		16#6636# => X"00000000",
		16#6637# => X"00000000",
		16#6638# => X"00000000",
		16#6639# => X"00000000",
		16#663a# => X"00000000",
		16#663b# => X"00000000",
		16#663c# => X"00000000",
		16#663d# => X"00000000",
		16#663e# => X"00000000",
		16#663f# => X"00000000",
		16#6640# => X"00000000",
		16#6641# => X"00000000",
		16#6642# => X"00000000",
		16#6643# => X"00000000",
		16#6644# => X"00000000",
		16#6645# => X"00000000",
		16#6646# => X"00000000",
		16#6647# => X"00000000",
		16#6648# => X"00000000",
		16#6649# => X"00000000",
		16#664a# => X"00000000",
		16#664b# => X"00000000",
		16#664c# => X"00000000",
		16#664d# => X"00000000",
		16#664e# => X"00000000",
		16#664f# => X"00000000",
		16#6650# => X"00000000",
		16#6651# => X"00000000",
		16#6652# => X"00000000",
		16#6653# => X"00000000",
		16#6654# => X"00000000",
		16#6655# => X"00000000",
		16#6656# => X"00000000",
		16#6657# => X"00000000",
		16#6658# => X"00000000",
		16#6659# => X"00000000",
		16#665a# => X"00000000",
		16#665b# => X"00000000",
		16#665c# => X"00000000",
		16#665d# => X"00000000",
		16#665e# => X"00000000",
		16#665f# => X"00000000",
		16#6660# => X"00000000",
		16#6661# => X"00000000",
		16#6662# => X"00000000",
		16#6663# => X"00000000",
		16#6664# => X"00000000",
		16#6665# => X"00000000",
		16#6666# => X"00000000",
		16#6667# => X"00000000",
		16#6668# => X"00000000",
		16#6669# => X"00000000",
		16#666a# => X"00000000",
		16#666b# => X"00000000",
		16#666c# => X"00000000",
		16#666d# => X"00000000",
		16#666e# => X"00000000",
		16#666f# => X"00000000",
		16#6670# => X"00000000",
		16#6671# => X"00000000",
		16#6672# => X"00000000",
		16#6673# => X"00000000",
		16#6674# => X"00000000",
		16#6675# => X"00000000",
		16#6676# => X"00000000",
		16#6677# => X"00000000",
		16#6678# => X"00000000",
		16#6679# => X"00000000",
		16#667a# => X"00000000",
		16#667b# => X"00000000",
		16#667c# => X"00000000",
		16#667d# => X"00000000",
		16#667e# => X"00000000",
		16#667f# => X"00000000",
		16#6680# => X"00000000",
		16#6681# => X"00000000",
		16#6682# => X"00000000",
		16#6683# => X"00000000",
		16#6684# => X"00000000",
		16#6685# => X"00000000",
		16#6686# => X"00000000",
		16#6687# => X"00000000",
		16#6688# => X"00000000",
		16#6689# => X"00000000",
		16#668a# => X"00000000",
		16#668b# => X"00000000",
		16#668c# => X"00000000",
		16#668d# => X"00000000",
		16#668e# => X"00000000",
		16#668f# => X"00000000",
		16#6690# => X"00000000",
		16#6691# => X"00000000",
		16#6692# => X"00000000",
		16#6693# => X"00000000",
		16#6694# => X"00000000",
		16#6695# => X"00000000",
		16#6696# => X"00000000",
		16#6697# => X"00000000",
		16#6698# => X"00000000",
		16#6699# => X"00000000",
		16#669a# => X"00000000",
		16#669b# => X"00000000",
		16#669c# => X"00000000",
		16#669d# => X"00000000",
		16#669e# => X"00000000",
		16#669f# => X"00000000",
		16#66a0# => X"00000000",
		16#66a1# => X"00000000",
		16#66a2# => X"00000000",
		16#66a3# => X"00000000",
		16#66a4# => X"00000000",
		16#66a5# => X"00000000",
		16#66a6# => X"00000000",
		16#66a7# => X"00000000",
		16#66a8# => X"00000000",
		16#66a9# => X"00000000",
		16#66aa# => X"00000000",
		16#66ab# => X"00000000",
		16#66ac# => X"00000000",
		16#66ad# => X"00000000",
		16#66ae# => X"00000000",
		16#66af# => X"00000000",
		16#66b0# => X"00000000",
		16#66b1# => X"00000000",
		16#66b2# => X"00000000",
		16#66b3# => X"00000000",
		16#66b4# => X"00000000",
		16#66b5# => X"00000000",
		16#66b6# => X"00000000",
		16#66b7# => X"00000000",
		16#66b8# => X"00000000",
		16#66b9# => X"00000000",
		16#66ba# => X"00000000",
		16#66bb# => X"00000000",
		16#66bc# => X"00000000",
		16#66bd# => X"00000000",
		16#66be# => X"00000000",
		16#66bf# => X"00000000",
		16#66c0# => X"00000000",
		16#66c1# => X"00000000",
		16#66c2# => X"00000000",
		16#66c3# => X"00000000",
		16#66c4# => X"00000000",
		16#66c5# => X"00000000",
		16#66c6# => X"00000000",
		16#66c7# => X"00000000",
		16#66c8# => X"00000000",
		16#66c9# => X"00000000",
		16#66ca# => X"00000000",
		16#66cb# => X"00000000",
		16#66cc# => X"00000000",
		16#66cd# => X"00000000",
		16#66ce# => X"00000000",
		16#66cf# => X"00000000",
		16#66d0# => X"00000000",
		16#66d1# => X"00000000",
		16#66d2# => X"00000000",
		16#66d3# => X"00000000",
		16#66d4# => X"00000000",
		16#66d5# => X"00000000",
		16#66d6# => X"00000000",
		16#66d7# => X"00000000",
		16#66d8# => X"00000000",
		16#66d9# => X"00000000",
		16#66da# => X"00000000",
		16#66db# => X"00000000",
		16#66dc# => X"00000000",
		16#66dd# => X"00000000",
		16#66de# => X"00000000",
		16#66df# => X"00000000",
		16#66e0# => X"00000000",
		16#66e1# => X"00000000",
		16#66e2# => X"00000000",
		16#66e3# => X"00000000",
		16#66e4# => X"00000000",
		16#66e5# => X"00000000",
		16#66e6# => X"00000000",
		16#66e7# => X"00000000",
		16#66e8# => X"00000000",
		16#66e9# => X"00000000",
		16#66ea# => X"00000000",
		16#66eb# => X"00000000",
		16#66ec# => X"00000000",
		16#66ed# => X"00000000",
		16#66ee# => X"00000000",
		16#66ef# => X"00000000",
		16#66f0# => X"00000000",
		16#66f1# => X"00000000",
		16#66f2# => X"00000000",
		16#66f3# => X"00000000",
		16#66f4# => X"00000000",
		16#66f5# => X"00000000",
		16#66f6# => X"00000000",
		16#66f7# => X"00000000",
		16#66f8# => X"00000000",
		16#66f9# => X"00000000",
		16#66fa# => X"00000000",
		16#66fb# => X"00000000",
		16#66fc# => X"00000000",
		16#66fd# => X"00000000",
		16#66fe# => X"00000000",
		16#66ff# => X"00000000",
		16#6700# => X"00000000",
		16#6701# => X"00000000",
		16#6702# => X"00000000",
		16#6703# => X"00000000",
		16#6704# => X"00000000",
		16#6705# => X"00000000",
		16#6706# => X"00000000",
		16#6707# => X"00000000",
		16#6708# => X"00000000",
		16#6709# => X"00000000",
		16#670a# => X"00000000",
		16#670b# => X"00000000",
		16#670c# => X"00000000",
		16#670d# => X"00000000",
		16#670e# => X"00000000",
		16#670f# => X"00000000",
		16#6710# => X"00000000",
		16#6711# => X"00000000",
		16#6712# => X"00000000",
		16#6713# => X"00000000",
		16#6714# => X"00000000",
		16#6715# => X"00000000",
		16#6716# => X"00000000",
		16#6717# => X"00000000",
		16#6718# => X"00000000",
		16#6719# => X"00000000",
		16#671a# => X"00000000",
		16#671b# => X"00000000",
		16#671c# => X"00000000",
		16#671d# => X"00000000",
		16#671e# => X"00000000",
		16#671f# => X"00000000",
		16#6720# => X"00000000",
		16#6721# => X"00000000",
		16#6722# => X"00000000",
		16#6723# => X"00000000",
		16#6724# => X"00000000",
		16#6725# => X"00000000",
		16#6726# => X"00000000",
		16#6727# => X"00000000",
		16#6728# => X"00000000",
		16#6729# => X"00000000",
		16#672a# => X"00000000",
		16#672b# => X"00000000",
		16#672c# => X"00000000",
		16#672d# => X"00000000",
		16#672e# => X"00000000",
		16#672f# => X"00000000",
		16#6730# => X"00000000",
		16#6731# => X"00000000",
		16#6732# => X"00000000",
		16#6733# => X"00000000",
		16#6734# => X"00000000",
		16#6735# => X"00000000",
		16#6736# => X"00000000",
		16#6737# => X"00000000",
		16#6738# => X"00000000",
		16#6739# => X"00000000",
		16#673a# => X"00000000",
		16#673b# => X"00000000",
		16#673c# => X"00000000",
		16#673d# => X"00000000",
		16#673e# => X"00000000",
		16#673f# => X"00000000",
		16#6740# => X"00000000",
		16#6741# => X"00000000",
		16#6742# => X"00000000",
		16#6743# => X"00000000",
		16#6744# => X"00000000",
		16#6745# => X"00000000",
		16#6746# => X"00000000",
		16#6747# => X"00000000",
		16#6748# => X"00000000",
		16#6749# => X"00000000",
		16#674a# => X"00000000",
		16#674b# => X"00000000",
		16#674c# => X"00000000",
		16#674d# => X"00000000",
		16#674e# => X"00000000",
		16#674f# => X"00000000",
		16#6750# => X"00000000",
		16#6751# => X"00000000",
		16#6752# => X"00000000",
		16#6753# => X"00000000",
		16#6754# => X"00000000",
		16#6755# => X"00000000",
		16#6756# => X"00000000",
		16#6757# => X"00000000",
		16#6758# => X"00000000",
		16#6759# => X"00000000",
		16#675a# => X"00000000",
		16#675b# => X"00000000",
		16#675c# => X"00000000",
		16#675d# => X"00000000",
		16#675e# => X"00000000",
		16#675f# => X"00000000",
		16#6760# => X"00000000",
		16#6761# => X"00000000",
		16#6762# => X"00000000",
		16#6763# => X"00000000",
		16#6764# => X"00000000",
		16#6765# => X"00000000",
		16#6766# => X"00000000",
		16#6767# => X"00000000",
		16#6768# => X"00000000",
		16#6769# => X"00000000",
		16#676a# => X"00000000",
		16#676b# => X"00000000",
		16#676c# => X"00000000",
		16#676d# => X"00000000",
		16#676e# => X"00000000",
		16#676f# => X"00000000",
		16#6770# => X"00000000",
		16#6771# => X"00000000",
		16#6772# => X"00000000",
		16#6773# => X"00000000",
		16#6774# => X"00000000",
		16#6775# => X"00000000",
		16#6776# => X"00000000",
		16#6777# => X"00000000",
		16#6778# => X"00000000",
		16#6779# => X"00000000",
		16#677a# => X"00000000",
		16#677b# => X"00000000",
		16#677c# => X"00000000",
		16#677d# => X"00000000",
		16#677e# => X"00000000",
		16#677f# => X"00000000",
		16#6780# => X"00000000",
		16#6781# => X"00000000",
		16#6782# => X"00000000",
		16#6783# => X"00000000",
		16#6784# => X"00000000",
		16#6785# => X"00000000",
		16#6786# => X"00000000",
		16#6787# => X"00000000",
		16#6788# => X"00000000",
		16#6789# => X"00000000",
		16#678a# => X"00000000",
		16#678b# => X"00000000",
		16#678c# => X"00000000",
		16#678d# => X"00000000",
		16#678e# => X"00000000",
		16#678f# => X"00000000",
		16#6790# => X"00000000",
		16#6791# => X"00000000",
		16#6792# => X"00000000",
		16#6793# => X"00000000",
		16#6794# => X"00000000",
		16#6795# => X"00000000",
		16#6796# => X"00000000",
		16#6797# => X"00000000",
		16#6798# => X"00000000",
		16#6799# => X"00000000",
		16#679a# => X"00000000",
		16#679b# => X"00000000",
		16#679c# => X"00000000",
		16#679d# => X"00000000",
		16#679e# => X"00000000",
		16#679f# => X"00000000",
		16#67a0# => X"00000000",
		16#67a1# => X"00000000",
		16#67a2# => X"00000000",
		16#67a3# => X"00000000",
		16#67a4# => X"00000000",
		16#67a5# => X"00000000",
		16#67a6# => X"00000000",
		16#67a7# => X"00000000",
		16#67a8# => X"00000000",
		16#67a9# => X"00000000",
		16#67aa# => X"00000000",
		16#67ab# => X"00000000",
		16#67ac# => X"00000000",
		16#67ad# => X"00000000",
		16#67ae# => X"00000000",
		16#67af# => X"00000000",
		16#67b0# => X"00000000",
		16#67b1# => X"00000000",
		16#67b2# => X"00000000",
		16#67b3# => X"00000000",
		16#67b4# => X"00000000",
		16#67b5# => X"00000000",
		16#67b6# => X"00000000",
		16#67b7# => X"00000000",
		16#67b8# => X"00000000",
		16#67b9# => X"00000000",
		16#67ba# => X"00000000",
		16#67bb# => X"00000000",
		16#67bc# => X"00000000",
		16#67bd# => X"00000000",
		16#67be# => X"00000000",
		16#67bf# => X"00000000",
		16#67c0# => X"00000000",
		16#67c1# => X"00000000",
		16#67c2# => X"00000000",
		16#67c3# => X"00000000",
		16#67c4# => X"00000000",
		16#67c5# => X"00000000",
		16#67c6# => X"00000000",
		16#67c7# => X"00000000",
		16#67c8# => X"00000000",
		16#67c9# => X"00000000",
		16#67ca# => X"00000000",
		16#67cb# => X"00000000",
		16#67cc# => X"00000000",
		16#67cd# => X"00000000",
		16#67ce# => X"00000000",
		16#67cf# => X"00000000",
		16#67d0# => X"00000000",
		16#67d1# => X"00000000",
		16#67d2# => X"00000000",
		16#67d3# => X"00000000",
		16#67d4# => X"00000000",
		16#67d5# => X"00000000",
		16#67d6# => X"00000000",
		16#67d7# => X"00000000",
		16#67d8# => X"00000000",
		16#67d9# => X"00000000",
		16#67da# => X"00000000",
		16#67db# => X"00000000",
		16#67dc# => X"00000000",
		16#67dd# => X"00000000",
		16#67de# => X"00000000",
		16#67df# => X"00000000",
		16#67e0# => X"00000000",
		16#67e1# => X"00000000",
		16#67e2# => X"00000000",
		16#67e3# => X"00000000",
		16#67e4# => X"00000000",
		16#67e5# => X"00000000",
		16#67e6# => X"00000000",
		16#67e7# => X"00000000",
		16#67e8# => X"00000000",
		16#67e9# => X"00000000",
		16#67ea# => X"00000000",
		16#67eb# => X"00000000",
		16#67ec# => X"00000000",
		16#67ed# => X"00000000",
		16#67ee# => X"00000000",
		16#67ef# => X"00000000",
		16#67f0# => X"00000000",
		16#67f1# => X"00000000",
		16#67f2# => X"00000000",
		16#67f3# => X"00000000",
		16#67f4# => X"00000000",
		16#67f5# => X"00000000",
		16#67f6# => X"00000000",
		16#67f7# => X"00000000",
		16#67f8# => X"00000000",
		16#67f9# => X"00000000",
		16#67fa# => X"00000000",
		16#67fb# => X"00000000",
		16#67fc# => X"00000000",
		16#67fd# => X"00000000",
		16#67fe# => X"00000000",
		16#67ff# => X"00000000",
		16#6800# => X"00000000",
		16#6801# => X"00000000",
		16#6802# => X"00000000",
		16#6803# => X"00000000",
		16#6804# => X"00000000",
		16#6805# => X"00000000",
		16#6806# => X"00000000",
		16#6807# => X"00000000",
		16#6808# => X"00000000",
		16#6809# => X"00000000",
		16#680a# => X"00000000",
		16#680b# => X"00000000",
		16#680c# => X"00000000",
		16#680d# => X"00000000",
		16#680e# => X"00000000",
		16#680f# => X"00000000",
		16#6810# => X"00000000",
		16#6811# => X"00000000",
		16#6812# => X"00000000",
		16#6813# => X"00000000",
		16#6814# => X"00000000",
		16#6815# => X"00000000",
		16#6816# => X"00000000",
		16#6817# => X"00000000",
		16#6818# => X"00000000",
		16#6819# => X"00000000",
		16#681a# => X"00000000",
		16#681b# => X"00000000",
		16#681c# => X"00000000",
		16#681d# => X"00000000",
		16#681e# => X"00000000",
		16#681f# => X"00000000",
		16#6820# => X"00000000",
		16#6821# => X"00000000",
		16#6822# => X"00000000",
		16#6823# => X"00000000",
		16#6824# => X"00000000",
		16#6825# => X"00000000",
		16#6826# => X"00000000",
		16#6827# => X"00000000",
		16#6828# => X"00000000",
		16#6829# => X"00000000",
		16#682a# => X"00000000",
		16#682b# => X"00000000",
		16#682c# => X"00000000",
		16#682d# => X"00000000",
		16#682e# => X"00000000",
		16#682f# => X"00000000",
		16#6830# => X"00000000",
		16#6831# => X"00000000",
		16#6832# => X"00000000",
		16#6833# => X"00000000",
		16#6834# => X"00000000",
		16#6835# => X"00000000",
		16#6836# => X"00000000",
		16#6837# => X"00000000",
		16#6838# => X"00000000",
		16#6839# => X"00000000",
		16#683a# => X"00000000",
		16#683b# => X"00000000",
		16#683c# => X"00000000",
		16#683d# => X"00000000",
		16#683e# => X"00000000",
		16#683f# => X"00000000",
		16#6840# => X"00000000",
		16#6841# => X"00000000",
		16#6842# => X"00000000",
		16#6843# => X"00000000",
		16#6844# => X"00000000",
		16#6845# => X"00000000",
		16#6846# => X"00000000",
		16#6847# => X"00000000",
		16#6848# => X"00000000",
		16#6849# => X"00000000",
		16#684a# => X"00000000",
		16#684b# => X"00000000",
		16#684c# => X"00000000",
		16#684d# => X"00000000",
		16#684e# => X"00000000",
		16#684f# => X"00000000",
		16#6850# => X"00000000",
		16#6851# => X"00000000",
		16#6852# => X"00000000",
		16#6853# => X"00000000",
		16#6854# => X"00000000",
		16#6855# => X"00000000",
		16#6856# => X"00000000",
		16#6857# => X"00000000",
		16#6858# => X"00000000",
		16#6859# => X"00000000",
		16#685a# => X"00000000",
		16#685b# => X"00000000",
		16#685c# => X"00000000",
		16#685d# => X"00000000",
		16#685e# => X"00000000",
		16#685f# => X"00000000",
		16#6860# => X"00000000",
		16#6861# => X"00000000",
		16#6862# => X"00000000",
		16#6863# => X"00000000",
		16#6864# => X"00000000",
		16#6865# => X"00000000",
		16#6866# => X"00000000",
		16#6867# => X"00000000",
		16#6868# => X"00000000",
		16#6869# => X"00000000",
		16#686a# => X"00000000",
		16#686b# => X"00000000",
		16#686c# => X"00000000",
		16#686d# => X"00000000",
		16#686e# => X"00000000",
		16#686f# => X"00000000",
		16#6870# => X"00000000",
		16#6871# => X"00000000",
		16#6872# => X"00000000",
		16#6873# => X"00000000",
		16#6874# => X"00000000",
		16#6875# => X"00000000",
		16#6876# => X"00000000",
		16#6877# => X"00000000",
		16#6878# => X"00000000",
		16#6879# => X"00000000",
		16#687a# => X"00000000",
		16#687b# => X"00000000",
		16#687c# => X"00000000",
		16#687d# => X"00000000",
		16#687e# => X"00000000",
		16#687f# => X"00000000",
		16#6880# => X"00000000",
		16#6881# => X"00000000",
		16#6882# => X"00000000",
		16#6883# => X"00000000",
		16#6884# => X"00000000",
		16#6885# => X"00000000",
		16#6886# => X"00000000",
		16#6887# => X"00000000",
		16#6888# => X"00000000",
		16#6889# => X"00000000",
		16#688a# => X"00000000",
		16#688b# => X"00000000",
		16#688c# => X"00000000",
		16#688d# => X"00000000",
		16#688e# => X"00000000",
		16#688f# => X"00000000",
		16#6890# => X"00000000",
		16#6891# => X"00000000",
		16#6892# => X"00000000",
		16#6893# => X"00000000",
		16#6894# => X"00000000",
		16#6895# => X"00000000",
		16#6896# => X"00000000",
		16#6897# => X"00000000",
		16#6898# => X"00000000",
		16#6899# => X"00000000",
		16#689a# => X"00000000",
		16#689b# => X"00000000",
		16#689c# => X"00000000",
		16#689d# => X"00000000",
		16#689e# => X"00000000",
		16#689f# => X"00000000",
		16#68a0# => X"00000000",
		16#68a1# => X"00000000",
		16#68a2# => X"00000000",
		16#68a3# => X"00000000",
		16#68a4# => X"00000000",
		16#68a5# => X"00000000",
		16#68a6# => X"00000000",
		16#68a7# => X"00000000",
		16#68a8# => X"00000000",
		16#68a9# => X"00000000",
		16#68aa# => X"00000000",
		16#68ab# => X"00000000",
		16#68ac# => X"00000000",
		16#68ad# => X"00000000",
		16#68ae# => X"00000000",
		16#68af# => X"00000000",
		16#68b0# => X"00000000",
		16#68b1# => X"00000000",
		16#68b2# => X"00000000",
		16#68b3# => X"00000000",
		16#68b4# => X"00000000",
		16#68b5# => X"00000000",
		16#68b6# => X"00000000",
		16#68b7# => X"00000000",
		16#68b8# => X"00000000",
		16#68b9# => X"00000000",
		16#68ba# => X"00000000",
		16#68bb# => X"00000000",
		16#68bc# => X"00000000",
		16#68bd# => X"00000000",
		16#68be# => X"00000000",
		16#68bf# => X"00000000",
		16#68c0# => X"00000000",
		16#68c1# => X"00000000",
		16#68c2# => X"00000000",
		16#68c3# => X"00000000",
		16#68c4# => X"00000000",
		16#68c5# => X"00000000",
		16#68c6# => X"00000000",
		16#68c7# => X"00000000",
		16#68c8# => X"00000000",
		16#68c9# => X"00000000",
		16#68ca# => X"00000000",
		16#68cb# => X"00000000",
		16#68cc# => X"00000000",
		16#68cd# => X"00000000",
		16#68ce# => X"00000000",
		16#68cf# => X"00000000",
		16#68d0# => X"00000000",
		16#68d1# => X"00000000",
		16#68d2# => X"00000000",
		16#68d3# => X"00000000",
		16#68d4# => X"00000000",
		16#68d5# => X"00000000",
		16#68d6# => X"00000000",
		16#68d7# => X"00000000",
		16#68d8# => X"00000000",
		16#68d9# => X"00000000",
		16#68da# => X"00000000",
		16#68db# => X"00000000",
		16#68dc# => X"00000000",
		16#68dd# => X"00000000",
		16#68de# => X"00000000",
		16#68df# => X"00000000",
		16#68e0# => X"00000000",
		16#68e1# => X"00000000",
		16#68e2# => X"00000000",
		16#68e3# => X"00000000",
		16#68e4# => X"00000000",
		16#68e5# => X"00000000",
		16#68e6# => X"00000000",
		16#68e7# => X"00000000",
		16#68e8# => X"00000000",
		16#68e9# => X"00000000",
		16#68ea# => X"00000000",
		16#68eb# => X"00000000",
		16#68ec# => X"00000000",
		16#68ed# => X"00000000",
		16#68ee# => X"00000000",
		16#68ef# => X"00000000",
		16#68f0# => X"00000000",
		16#68f1# => X"00000000",
		16#68f2# => X"00000000",
		16#68f3# => X"00000000",
		16#68f4# => X"00000000",
		16#68f5# => X"00000000",
		16#68f6# => X"00000000",
		16#68f7# => X"00000000",
		16#68f8# => X"00000000",
		16#68f9# => X"00000000",
		16#68fa# => X"00000000",
		16#68fb# => X"00000000",
		16#68fc# => X"00000000",
		16#68fd# => X"00000000",
		16#68fe# => X"00000000",
		16#68ff# => X"00000000",
		16#6900# => X"00000000",
		16#6901# => X"00000000",
		16#6902# => X"00000000",
		16#6903# => X"00000000",
		16#6904# => X"00000000",
		16#6905# => X"00000000",
		16#6906# => X"00000000",
		16#6907# => X"00000000",
		16#6908# => X"00000000",
		16#6909# => X"00000000",
		16#690a# => X"00000000",
		16#690b# => X"00000000",
		16#690c# => X"00000000",
		16#690d# => X"00000000",
		16#690e# => X"00000000",
		16#690f# => X"00000000",
		16#6910# => X"00000000",
		16#6911# => X"00000000",
		16#6912# => X"00000000",
		16#6913# => X"00000000",
		16#6914# => X"00000000",
		16#6915# => X"00000000",
		16#6916# => X"00000000",
		16#6917# => X"00000000",
		16#6918# => X"00000000",
		16#6919# => X"00000000",
		16#691a# => X"00000000",
		16#691b# => X"00000000",
		16#691c# => X"00000000",
		16#691d# => X"00000000",
		16#691e# => X"00000000",
		16#691f# => X"00000000",
		16#6920# => X"00000000",
		16#6921# => X"00000000",
		16#6922# => X"00000000",
		16#6923# => X"00000000",
		16#6924# => X"00000000",
		16#6925# => X"00000000",
		16#6926# => X"00000000",
		16#6927# => X"00000000",
		16#6928# => X"00000000",
		16#6929# => X"00000000",
		16#692a# => X"00000000",
		16#692b# => X"00000000",
		16#692c# => X"00000000",
		16#692d# => X"00000000",
		16#692e# => X"00000000",
		16#692f# => X"00000000",
		16#6930# => X"00000000",
		16#6931# => X"00000000",
		16#6932# => X"00000000",
		16#6933# => X"00000000",
		16#6934# => X"00000000",
		16#6935# => X"00000000",
		16#6936# => X"00000000",
		16#6937# => X"00000000",
		16#6938# => X"00000000",
		16#6939# => X"00000000",
		16#693a# => X"00000000",
		16#693b# => X"00000000",
		16#693c# => X"00000000",
		16#693d# => X"00000000",
		16#693e# => X"00000000",
		16#693f# => X"00000000",
		16#6940# => X"00000000",
		16#6941# => X"00000000",
		16#6942# => X"00000000",
		16#6943# => X"00000000",
		16#6944# => X"00000000",
		16#6945# => X"00000000",
		16#6946# => X"00000000",
		16#6947# => X"00000000",
		16#6948# => X"00000000",
		16#6949# => X"00000000",
		16#694a# => X"00000000",
		16#694b# => X"00000000",
		16#694c# => X"00000000",
		16#694d# => X"00000000",
		16#694e# => X"00000000",
		16#694f# => X"00000000",
		16#6950# => X"00000000",
		16#6951# => X"00000000",
		16#6952# => X"00000000",
		16#6953# => X"00000000",
		16#6954# => X"00000000",
		16#6955# => X"00000000",
		16#6956# => X"00000000",
		16#6957# => X"00000000",
		16#6958# => X"00000000",
		16#6959# => X"00000000",
		16#695a# => X"00000000",
		16#695b# => X"00000000",
		16#695c# => X"00000000",
		16#695d# => X"00000000",
		16#695e# => X"00000000",
		16#695f# => X"00000000",
		16#6960# => X"00000000",
		16#6961# => X"00000000",
		16#6962# => X"00000000",
		16#6963# => X"00000000",
		16#6964# => X"00000000",
		16#6965# => X"00000000",
		16#6966# => X"00000000",
		16#6967# => X"00000000",
		16#6968# => X"00000000",
		16#6969# => X"00000000",
		16#696a# => X"00000000",
		16#696b# => X"00000000",
		16#696c# => X"00000000",
		16#696d# => X"00000000",
		16#696e# => X"00000000",
		16#696f# => X"00000000",
		16#6970# => X"00000000",
		16#6971# => X"00000000",
		16#6972# => X"00000000",
		16#6973# => X"00000000",
		16#6974# => X"00000000",
		16#6975# => X"00000000",
		16#6976# => X"00000000",
		16#6977# => X"00000000",
		16#6978# => X"00000000",
		16#6979# => X"00000000",
		16#697a# => X"00000000",
		16#697b# => X"00000000",
		16#697c# => X"00000000",
		16#697d# => X"00000000",
		16#697e# => X"00000000",
		16#697f# => X"00000000",
		16#6980# => X"00000000",
		16#6981# => X"00000000",
		16#6982# => X"00000000",
		16#6983# => X"00000000",
		16#6984# => X"00000000",
		16#6985# => X"00000000",
		16#6986# => X"00000000",
		16#6987# => X"00000000",
		16#6988# => X"00000000",
		16#6989# => X"00000000",
		16#698a# => X"00000000",
		16#698b# => X"00000000",
		16#698c# => X"00000000",
		16#698d# => X"00000000",
		16#698e# => X"00000000",
		16#698f# => X"00000000",
		16#6990# => X"00000000",
		16#6991# => X"00000000",
		16#6992# => X"00000000",
		16#6993# => X"00000000",
		16#6994# => X"00000000",
		16#6995# => X"00000000",
		16#6996# => X"00000000",
		16#6997# => X"00000000",
		16#6998# => X"00000000",
		16#6999# => X"00000000",
		16#699a# => X"00000000",
		16#699b# => X"00000000",
		16#699c# => X"00000000",
		16#699d# => X"00000000",
		16#699e# => X"00000000",
		16#699f# => X"00000000",
		16#69a0# => X"00000000",
		16#69a1# => X"00000000",
		16#69a2# => X"00000000",
		16#69a3# => X"00000000",
		16#69a4# => X"00000000",
		16#69a5# => X"00000000",
		16#69a6# => X"00000000",
		16#69a7# => X"00000000",
		16#69a8# => X"00000000",
		16#69a9# => X"00000000",
		16#69aa# => X"00000000",
		16#69ab# => X"00000000",
		16#69ac# => X"00000000",
		16#69ad# => X"00000000",
		16#69ae# => X"00000000",
		16#69af# => X"00000000",
		16#69b0# => X"00000000",
		16#69b1# => X"00000000",
		16#69b2# => X"00000000",
		16#69b3# => X"00000000",
		16#69b4# => X"00000000",
		16#69b5# => X"00000000",
		16#69b6# => X"00000000",
		16#69b7# => X"00000000",
		16#69b8# => X"00000000",
		16#69b9# => X"00000000",
		16#69ba# => X"00000000",
		16#69bb# => X"00000000",
		16#69bc# => X"00000000",
		16#69bd# => X"00000000",
		16#69be# => X"00000000",
		16#69bf# => X"00000000",
		16#69c0# => X"00000000",
		16#69c1# => X"00000000",
		16#69c2# => X"00000000",
		16#69c3# => X"00000000",
		16#69c4# => X"00000000",
		16#69c5# => X"00000000",
		16#69c6# => X"00000000",
		16#69c7# => X"00000000",
		16#69c8# => X"00000000",
		16#69c9# => X"00000000",
		16#69ca# => X"00000000",
		16#69cb# => X"00000000",
		16#69cc# => X"00000000",
		16#69cd# => X"00000000",
		16#69ce# => X"00000000",
		16#69cf# => X"00000000",
		16#69d0# => X"00000000",
		16#69d1# => X"00000000",
		16#69d2# => X"00000000",
		16#69d3# => X"00000000",
		16#69d4# => X"00000000",
		16#69d5# => X"00000000",
		16#69d6# => X"00000000",
		16#69d7# => X"00000000",
		16#69d8# => X"00000000",
		16#69d9# => X"00000000",
		16#69da# => X"00000000",
		16#69db# => X"00000000",
		16#69dc# => X"00000000",
		16#69dd# => X"00000000",
		16#69de# => X"00000000",
		16#69df# => X"00000000",
		16#69e0# => X"00000000",
		16#69e1# => X"00000000",
		16#69e2# => X"00000000",
		16#69e3# => X"00000000",
		16#69e4# => X"00000000",
		16#69e5# => X"00000000",
		16#69e6# => X"00000000",
		16#69e7# => X"00000000",
		16#69e8# => X"00000000",
		16#69e9# => X"00000000",
		16#69ea# => X"00000000",
		16#69eb# => X"00000000",
		16#69ec# => X"00000000",
		16#69ed# => X"00000000",
		16#69ee# => X"00000000",
		16#69ef# => X"00000000",
		16#69f0# => X"00000000",
		16#69f1# => X"00000000",
		16#69f2# => X"00000000",
		16#69f3# => X"00000000",
		16#69f4# => X"00000000",
		16#69f5# => X"00000000",
		16#69f6# => X"00000000",
		16#69f7# => X"00000000",
		16#69f8# => X"00000000",
		16#69f9# => X"00000000",
		16#69fa# => X"00000000",
		16#69fb# => X"00000000",
		16#69fc# => X"00000000",
		16#69fd# => X"00000000",
		16#69fe# => X"00000000",
		16#69ff# => X"00000000",
		16#6a00# => X"00000000",
		16#6a01# => X"00000000",
		16#6a02# => X"00000000",
		16#6a03# => X"00000000",
		16#6a04# => X"00000000",
		16#6a05# => X"00000000",
		16#6a06# => X"00000000",
		16#6a07# => X"00000000",
		16#6a08# => X"00000000",
		16#6a09# => X"00000000",
		16#6a0a# => X"00000000",
		16#6a0b# => X"00000000",
		16#6a0c# => X"00000000",
		16#6a0d# => X"00000000",
		16#6a0e# => X"00000000",
		16#6a0f# => X"00000000",
		16#6a10# => X"00000000",
		16#6a11# => X"00000000",
		16#6a12# => X"00000000",
		16#6a13# => X"00000000",
		16#6a14# => X"00000000",
		16#6a15# => X"00000000",
		16#6a16# => X"00000000",
		16#6a17# => X"00000000",
		16#6a18# => X"00000000",
		16#6a19# => X"00000000",
		16#6a1a# => X"00000000",
		16#6a1b# => X"00000000",
		16#6a1c# => X"00000000",
		16#6a1d# => X"00000000",
		16#6a1e# => X"00000000",
		16#6a1f# => X"00000000",
		16#6a20# => X"00000000",
		16#6a21# => X"00000000",
		16#6a22# => X"00000000",
		16#6a23# => X"00000000",
		16#6a24# => X"00000000",
		16#6a25# => X"00000000",
		16#6a26# => X"00000000",
		16#6a27# => X"00000000",
		16#6a28# => X"00000000",
		16#6a29# => X"00000000",
		16#6a2a# => X"00000000",
		16#6a2b# => X"00000000",
		16#6a2c# => X"00000000",
		16#6a2d# => X"00000000",
		16#6a2e# => X"00000000",
		16#6a2f# => X"00000000",
		16#6a30# => X"00000000",
		16#6a31# => X"00000000",
		16#6a32# => X"00000000",
		16#6a33# => X"00000000",
		16#6a34# => X"00000000",
		16#6a35# => X"00000000",
		16#6a36# => X"00000000",
		16#6a37# => X"00000000",
		16#6a38# => X"00000000",
		16#6a39# => X"00000000",
		16#6a3a# => X"00000000",
		16#6a3b# => X"00000000",
		16#6a3c# => X"00000000",
		16#6a3d# => X"00000000",
		16#6a3e# => X"00000000",
		16#6a3f# => X"00000000",
		16#6a40# => X"00000000",
		16#6a41# => X"00000000",
		16#6a42# => X"00000000",
		16#6a43# => X"00000000",
		16#6a44# => X"00000000",
		16#6a45# => X"00000000",
		16#6a46# => X"00000000",
		16#6a47# => X"00000000",
		16#6a48# => X"00000000",
		16#6a49# => X"00000000",
		16#6a4a# => X"00000000",
		16#6a4b# => X"00000000",
		16#6a4c# => X"00000000",
		16#6a4d# => X"00000000",
		16#6a4e# => X"00000000",
		16#6a4f# => X"00000000",
		16#6a50# => X"00000000",
		16#6a51# => X"00000000",
		16#6a52# => X"00000000",
		16#6a53# => X"00000000",
		16#6a54# => X"00000000",
		16#6a55# => X"00000000",
		16#6a56# => X"00000000",
		16#6a57# => X"00000000",
		16#6a58# => X"00000000",
		16#6a59# => X"00000000",
		16#6a5a# => X"00000000",
		16#6a5b# => X"00000000",
		16#6a5c# => X"00000000",
		16#6a5d# => X"00000000",
		16#6a5e# => X"00000000",
		16#6a5f# => X"00000000",
		16#6a60# => X"00000000",
		16#6a61# => X"00000000",
		16#6a62# => X"00000000",
		16#6a63# => X"00000000",
		16#6a64# => X"00000000",
		16#6a65# => X"00000000",
		16#6a66# => X"00000000",
		16#6a67# => X"00000000",
		16#6a68# => X"00000000",
		16#6a69# => X"00000000",
		16#6a6a# => X"00000000",
		16#6a6b# => X"00000000",
		16#6a6c# => X"00000000",
		16#6a6d# => X"00000000",
		16#6a6e# => X"00000000",
		16#6a6f# => X"00000000",
		16#6a70# => X"00000000",
		16#6a71# => X"00000000",
		16#6a72# => X"00000000",
		16#6a73# => X"00000000",
		16#6a74# => X"00000000",
		16#6a75# => X"00000000",
		16#6a76# => X"00000000",
		16#6a77# => X"00000000",
		16#6a78# => X"00000000",
		16#6a79# => X"00000000",
		16#6a7a# => X"00000000",
		16#6a7b# => X"00000000",
		16#6a7c# => X"00000000",
		16#6a7d# => X"00000000",
		16#6a7e# => X"00000000",
		16#6a7f# => X"00000000",
		16#6a80# => X"00000000",
		16#6a81# => X"00000000",
		16#6a82# => X"00000000",
		16#6a83# => X"00000000",
		16#6a84# => X"00000000",
		16#6a85# => X"00000000",
		16#6a86# => X"00000000",
		16#6a87# => X"00000000",
		16#6a88# => X"00000000",
		16#6a89# => X"00000000",
		16#6a8a# => X"00000000",
		16#6a8b# => X"00000000",
		16#6a8c# => X"00000000",
		16#6a8d# => X"00000000",
		16#6a8e# => X"00000000",
		16#6a8f# => X"00000000",
		16#6a90# => X"00000000",
		16#6a91# => X"00000000",
		16#6a92# => X"00000000",
		16#6a93# => X"00000000",
		16#6a94# => X"00000000",
		16#6a95# => X"00000000",
		16#6a96# => X"00000000",
		16#6a97# => X"00000000",
		16#6a98# => X"00000000",
		16#6a99# => X"00000000",
		16#6a9a# => X"00000000",
		16#6a9b# => X"00000000",
		16#6a9c# => X"00000000",
		16#6a9d# => X"00000000",
		16#6a9e# => X"00000000",
		16#6a9f# => X"00000000",
		16#6aa0# => X"00000000",
		16#6aa1# => X"00000000",
		16#6aa2# => X"00000000",
		16#6aa3# => X"00000000",
		16#6aa4# => X"00000000",
		16#6aa5# => X"00000000",
		16#6aa6# => X"00000000",
		16#6aa7# => X"00000000",
		16#6aa8# => X"00000000",
		16#6aa9# => X"00000000",
		16#6aaa# => X"00000000",
		16#6aab# => X"00000000",
		16#6aac# => X"00000000",
		16#6aad# => X"00000000",
		16#6aae# => X"00000000",
		16#6aaf# => X"00000000",
		16#6ab0# => X"00000000",
		16#6ab1# => X"00000000",
		16#6ab2# => X"00000000",
		16#6ab3# => X"00000000",
		16#6ab4# => X"00000000",
		16#6ab5# => X"00000000",
		16#6ab6# => X"00000000",
		16#6ab7# => X"00000000",
		16#6ab8# => X"00000000",
		16#6ab9# => X"00000000",
		16#6aba# => X"00000000",
		16#6abb# => X"00000000",
		16#6abc# => X"00000000",
		16#6abd# => X"00000000",
		16#6abe# => X"00000000",
		16#6abf# => X"00000000",
		16#6ac0# => X"00000000",
		16#6ac1# => X"00000000",
		16#6ac2# => X"00000000",
		16#6ac3# => X"00000000",
		16#6ac4# => X"00000000",
		16#6ac5# => X"00000000",
		16#6ac6# => X"00000000",
		16#6ac7# => X"00000000",
		16#6ac8# => X"00000000",
		16#6ac9# => X"00000000",
		16#6aca# => X"00000000",
		16#6acb# => X"00000000",
		16#6acc# => X"00000000",
		16#6acd# => X"00000000",
		16#6ace# => X"00000000",
		16#6acf# => X"00000000",
		16#6ad0# => X"00000000",
		16#6ad1# => X"00000000",
		16#6ad2# => X"00000000",
		16#6ad3# => X"00000000",
		16#6ad4# => X"00000000",
		16#6ad5# => X"00000000",
		16#6ad6# => X"00000000",
		16#6ad7# => X"00000000",
		16#6ad8# => X"00000000",
		16#6ad9# => X"00000000",
		16#6ada# => X"00000000",
		16#6adb# => X"00000000",
		16#6adc# => X"00000000",
		16#6add# => X"00000000",
		16#6ade# => X"00000000",
		16#6adf# => X"00000000",
		16#6ae0# => X"00000000",
		16#6ae1# => X"00000000",
		16#6ae2# => X"00000000",
		16#6ae3# => X"00000000",
		16#6ae4# => X"00000000",
		16#6ae5# => X"00000000",
		16#6ae6# => X"00000000",
		16#6ae7# => X"00000000",
		16#6ae8# => X"00000000",
		16#6ae9# => X"00000000",
		16#6aea# => X"00000000",
		16#6aeb# => X"00000000",
		16#6aec# => X"00000000",
		16#6aed# => X"00000000",
		16#6aee# => X"00000000",
		16#6aef# => X"00000000",
		16#6af0# => X"00000000",
		16#6af1# => X"00000000",
		16#6af2# => X"00000000",
		16#6af3# => X"00000000",
		16#6af4# => X"00000000",
		16#6af5# => X"00000000",
		16#6af6# => X"00000000",
		16#6af7# => X"00000000",
		16#6af8# => X"00000000",
		16#6af9# => X"00000000",
		16#6afa# => X"00000000",
		16#6afb# => X"00000000",
		16#6afc# => X"00000000",
		16#6afd# => X"00000000",
		16#6afe# => X"00000000",
		16#6aff# => X"00000000",
		16#6b00# => X"00000000",
		16#6b01# => X"00000000",
		16#6b02# => X"00000000",
		16#6b03# => X"00000000",
		16#6b04# => X"00000000",
		16#6b05# => X"00000000",
		16#6b06# => X"00000000",
		16#6b07# => X"00000000",
		16#6b08# => X"00000000",
		16#6b09# => X"00000000",
		16#6b0a# => X"00000000",
		16#6b0b# => X"00000000",
		16#6b0c# => X"00000000",
		16#6b0d# => X"00000000",
		16#6b0e# => X"00000000",
		16#6b0f# => X"00000000",
		16#6b10# => X"00000000",
		16#6b11# => X"00000000",
		16#6b12# => X"00000000",
		16#6b13# => X"00000000",
		16#6b14# => X"00000000",
		16#6b15# => X"00000000",
		16#6b16# => X"00000000",
		16#6b17# => X"00000000",
		16#6b18# => X"00000000",
		16#6b19# => X"00000000",
		16#6b1a# => X"00000000",
		16#6b1b# => X"00000000",
		16#6b1c# => X"00000000",
		16#6b1d# => X"00000000",
		16#6b1e# => X"00000000",
		16#6b1f# => X"00000000",
		16#6b20# => X"00000000",
		16#6b21# => X"00000000",
		16#6b22# => X"00000000",
		16#6b23# => X"00000000",
		16#6b24# => X"00000000",
		16#6b25# => X"00000000",
		16#6b26# => X"00000000",
		16#6b27# => X"00000000",
		16#6b28# => X"00000000",
		16#6b29# => X"00000000",
		16#6b2a# => X"00000000",
		16#6b2b# => X"00000000",
		16#6b2c# => X"00000000",
		16#6b2d# => X"00000000",
		16#6b2e# => X"00000000",
		16#6b2f# => X"00000000",
		16#6b30# => X"00000000",
		16#6b31# => X"00000000",
		16#6b32# => X"00000000",
		16#6b33# => X"00000000",
		16#6b34# => X"00000000",
		16#6b35# => X"00000000",
		16#6b36# => X"00000000",
		16#6b37# => X"00000000",
		16#6b38# => X"00000000",
		16#6b39# => X"00000000",
		16#6b3a# => X"00000000",
		16#6b3b# => X"00000000",
		16#6b3c# => X"00000000",
		16#6b3d# => X"00000000",
		16#6b3e# => X"00000000",
		16#6b3f# => X"00000000",
		16#6b40# => X"00000000",
		16#6b41# => X"00000000",
		16#6b42# => X"00000000",
		16#6b43# => X"00000000",
		16#6b44# => X"00000000",
		16#6b45# => X"00000000",
		16#6b46# => X"00000000",
		16#6b47# => X"00000000",
		16#6b48# => X"00000000",
		16#6b49# => X"00000000",
		16#6b4a# => X"00000000",
		16#6b4b# => X"00000000",
		16#6b4c# => X"00000000",
		16#6b4d# => X"00000000",
		16#6b4e# => X"00000000",
		16#6b4f# => X"00000000",
		16#6b50# => X"00000000",
		16#6b51# => X"00000000",
		16#6b52# => X"00000000",
		16#6b53# => X"00000000",
		16#6b54# => X"00000000",
		16#6b55# => X"00000000",
		16#6b56# => X"00000000",
		16#6b57# => X"00000000",
		16#6b58# => X"00000000",
		16#6b59# => X"00000000",
		16#6b5a# => X"00000000",
		16#6b5b# => X"00000000",
		16#6b5c# => X"00000000",
		16#6b5d# => X"00000000",
		16#6b5e# => X"00000000",
		16#6b5f# => X"00000000",
		16#6b60# => X"00000000",
		16#6b61# => X"00000000",
		16#6b62# => X"00000000",
		16#6b63# => X"00000000",
		16#6b64# => X"00000000",
		16#6b65# => X"00000000",
		16#6b66# => X"00000000",
		16#6b67# => X"00000000",
		16#6b68# => X"00000000",
		16#6b69# => X"00000000",
		16#6b6a# => X"00000000",
		16#6b6b# => X"00000000",
		16#6b6c# => X"ffffffff",
		16#6b6d# => X"00000000",
		16#6b6e# => X"ffffffff",
		16#6b6f# => X"00000000",
		16#6b70# => X"00000000",
		16#6b71# => X"00000000",
		16#6b72# => X"00000000",
		16#6b73# => X"0001834c",
		16#6b74# => X"00018353",
		16#6b75# => X"00018358",
		16#6b76# => X"00000066",
		16#6b77# => X"00000001",
		16#6b78# => X"00000008",
		16#6b79# => X"0001ade8",
		16#6b7a# => X"00000000",
		16#6b7b# => X"0001b0d4",
		16#6b7c# => X"0001b13c",
		16#6b7d# => X"0001b1a4",
		16#6b7e# => X"00000000",
		16#6b7f# => X"00000000",
		16#6b80# => X"00000000",
		16#6b81# => X"00000000",
		16#6b82# => X"00000000",
		16#6b83# => X"00000000",
		16#6b84# => X"00000000",
		16#6b85# => X"00000000",
		16#6b86# => X"00000000",
		16#6b87# => X"00018894",
		16#6b88# => X"00000000",
		16#6b89# => X"00000000",
		16#6b8a# => X"00000000",
		16#6b8b# => X"00000000",
		16#6b8c# => X"00000000",
		16#6b8d# => X"00000000",
		16#6b8e# => X"00000000",
		16#6b8f# => X"00000000",
		16#6b90# => X"00000000",
		16#6b91# => X"00000000",
		16#6b92# => X"00000000",
		16#6b93# => X"00000000",
		16#6b94# => X"00000000",
		16#6b95# => X"00000000",
		16#6b96# => X"00000000",
		16#6b97# => X"00000000",
		16#6b98# => X"00000000",
		16#6b99# => X"00000000",
		16#6b9a# => X"00000000",
		16#6b9b# => X"00000000",
		16#6b9c# => X"00000000",
		16#6b9d# => X"00000000",
		16#6b9e# => X"00000000",
		16#6b9f# => X"00000000",
		16#6ba0# => X"00000000",
		16#6ba1# => X"00000000",
		16#6ba2# => X"00000000",
		16#6ba3# => X"00000000",
		16#6ba4# => X"00000001",
		16#6ba5# => X"330eabcd",
		16#6ba6# => X"1234e66d",
		16#6ba7# => X"deec0005",
		16#6ba8# => X"000b0000",
		16#6ba9# => X"00000000",
		16#6baa# => X"00000000",
		16#6bab# => X"00000000",
		16#6bac# => X"00000000",
		16#6bad# => X"00000000",
		16#6bae# => X"00000000",
		16#6baf# => X"00000000",
		16#6bb0# => X"00000000",
		16#6bb1# => X"00000000",
		16#6bb2# => X"00000000",
		16#6bb3# => X"00000000",
		16#6bb4# => X"00000000",
		16#6bb5# => X"00000000",
		16#6bb6# => X"00000000",
		16#6bb7# => X"00000000",
		16#6bb8# => X"00000000",
		16#6bb9# => X"00000000",
		16#6bba# => X"00000000",
		16#6bbb# => X"00000000",
		16#6bbc# => X"00000000",
		16#6bbd# => X"00000000",
		16#6bbe# => X"00000000",
		16#6bbf# => X"00000000",
		16#6bc0# => X"00000000",
		16#6bc1# => X"00000000",
		16#6bc2# => X"00000000",
		16#6bc3# => X"00000000",
		16#6bc4# => X"00000000",
		16#6bc5# => X"00000000",
		16#6bc6# => X"00000000",
		16#6bc7# => X"00000000",
		16#6bc8# => X"00000000",
		16#6bc9# => X"00000000",
		16#6bca# => X"00000000",
		16#6bcb# => X"00000000",
		16#6bcc# => X"00000000",
		16#6bcd# => X"00000000",
		16#6bce# => X"00000000",
		16#6bcf# => X"00000000",
		16#6bd0# => X"00000000",
		16#6bd1# => X"00000000",
		16#6bd2# => X"00000000",
		16#6bd3# => X"00000000",
		16#6bd4# => X"00000000",
		16#6bd5# => X"00000000",
		16#6bd6# => X"00000000",
		16#6bd7# => X"00000000",
		16#6bd8# => X"00000000",
		16#6bd9# => X"00000000",
		16#6bda# => X"00000000",
		16#6bdb# => X"00000000",
		16#6bdc# => X"00000000",
		16#6bdd# => X"00000000",
		16#6bde# => X"00000000",
		16#6bdf# => X"00000000",
		16#6be0# => X"00000000",
		16#6be1# => X"00000000",
		16#6be2# => X"00000000",
		16#6be3# => X"00000000",
		16#6be4# => X"00000000",
		16#6be5# => X"00000000",
		16#6be6# => X"00000000",
		16#6be7# => X"00000000",
		16#6be8# => X"00000000",
		16#6be9# => X"00000000",
		16#6bea# => X"00000000",
		16#6beb# => X"00000000",
		16#6bec# => X"00000000",
		16#6bed# => X"00000000",
		16#6bee# => X"00000000",
		16#6bef# => X"00000000",
		16#6bf0# => X"00000000",
		16#6bf1# => X"00000000",
		16#6bf2# => X"00000000",
		16#6bf3# => X"00000000",
		16#6bf4# => X"00000000",
		16#6bf5# => X"00000000",
		16#6bf6# => X"00000000",
		16#6bf7# => X"00000000",
		16#6bf8# => X"00000000",
		16#6bf9# => X"00000000",
		16#6bfa# => X"00000000",
		16#6bfb# => X"00000000",
		16#6bfc# => X"00000000",
		16#6bfd# => X"00000000",
		16#6bfe# => X"00000000",
		16#6bff# => X"00000000",
		16#6c00# => X"00000000",
		16#6c01# => X"00000000",
		16#6c02# => X"00000000",
		16#6c03# => X"00000000",
		16#6c04# => X"00000000",
		16#6c05# => X"00000000",
		16#6c06# => X"00000000",
		16#6c07# => X"00000000",
		16#6c08# => X"00000000",
		16#6c09# => X"00000000",
		16#6c0a# => X"00000000",
		16#6c0b# => X"00000000",
		16#6c0c# => X"00000000",
		16#6c0d# => X"00000000",
		16#6c0e# => X"00000000",
		16#6c0f# => X"00000000",
		16#6c10# => X"00000000",
		16#6c11# => X"00000000",
		16#6c12# => X"00000000",
		16#6c13# => X"00000000",
		16#6c14# => X"00000000",
		16#6c15# => X"00000000",
		16#6c16# => X"00000000",
		16#6c17# => X"00000000",
		16#6c18# => X"00000000",
		16#6c19# => X"00000000",
		16#6c1a# => X"00000000",
		16#6c1b# => X"00000000",
		16#6c1c# => X"00000000",
		16#6c1d# => X"00000000",
		16#6c1e# => X"00000000",
		16#6c1f# => X"00000000",
		16#6c20# => X"00000000",
		16#6c21# => X"00000000",
		16#6c22# => X"00000000",
		16#6c23# => X"00000000",
		16#6c24# => X"00000000",
		16#6c25# => X"00000000",
		16#6c26# => X"00000000",
		16#6c27# => X"00000000",
		16#6c28# => X"00000000",
		16#6c29# => X"00000000",
		16#6c2a# => X"00000000",
		16#6c2b# => X"00000000",
		16#6c2c# => X"00000000",
		16#6c2d# => X"00000000",
		16#6c2e# => X"00000000",
		16#6c2f# => X"00000000",
		16#6c30# => X"00000000",
		16#6c31# => X"00000000",
		16#6c32# => X"00000000",
		16#6c33# => X"00000000",
		16#6c34# => X"00000000",
		16#6c35# => X"00000000",
		16#6c36# => X"00000000",
		16#6c37# => X"00000000",
		16#6c38# => X"00000000",
		16#6c39# => X"00000000",
		16#6c3a# => X"00000000",
		16#6c3b# => X"00000000",
		16#6c3c# => X"00000000",
		16#6c3d# => X"00000000",
		16#6c3e# => X"00000000",
		16#6c3f# => X"00000000",
		16#6c40# => X"00000000",
		16#6c41# => X"00000000",
		16#6c42# => X"00000000",
		16#6c43# => X"00000000",
		16#6c44# => X"00000000",
		16#6c45# => X"00000000",
		16#6c46# => X"00000000",
		16#6c47# => X"00000000",
		16#6c48# => X"00000000",
		16#6c49# => X"00000000",
		16#6c4a# => X"00000000",
		16#6c4b# => X"00000000",
		16#6c4c# => X"00000000",
		16#6c4d# => X"00000000",
		16#6c4e# => X"00000000",
		16#6c4f# => X"00000000",
		16#6c50# => X"00000000",
		16#6c51# => X"00000000",
		16#6c52# => X"00000000",
		16#6c53# => X"00000000",
		16#6c54# => X"00000000",
		16#6c55# => X"00000000",
		16#6c56# => X"00000000",
		16#6c57# => X"00000000",
		16#6c58# => X"00000000",
		16#6c59# => X"00000000",
		16#6c5a# => X"00000000",
		16#6c5b# => X"00000000",
		16#6c5c# => X"00000000",
		16#6c5d# => X"00000000",
		16#6c5e# => X"00000000",
		16#6c5f# => X"00000000",
		16#6c60# => X"00000000",
		16#6c61# => X"00000000",
		16#6c62# => X"00000000",
		16#6c63# => X"00000000",
		16#6c64# => X"00000000",
		16#6c65# => X"00000000",
		16#6c66# => X"00000000",
		16#6c67# => X"00000000",
		16#6c68# => X"00000000",
		16#6c69# => X"00000000",
		16#6c6a# => X"00000000",
		16#6c6b# => X"00000000",
		16#6c6c# => X"00000000",
		16#6c6d# => X"00000000",
		16#6c6e# => X"00000000",
		16#6c6f# => X"00000000",
		16#6c70# => X"00000000",
		16#6c71# => X"00000000",
		16#6c72# => X"00000000",
		16#6c73# => X"00000000",
		16#6c74# => X"00000000",
		16#6c75# => X"00000000",
		16#6c76# => X"00000000",
		16#6c77# => X"00000000",
		16#6c78# => X"00000000",
		16#6c79# => X"00000000",
		16#6c7a# => X"00000000",
		16#6c7b# => X"00000000",
		16#6c7c# => X"00000000",
		16#6c7d# => X"00000000",
		16#6c7e# => X"00000000",
		16#6c7f# => X"00000000",
		16#6c80# => X"00000000",
		16#6c81# => X"00000000",
		16#6c82# => X"00000000",
		16#6c83# => X"00000000",
		16#6c84# => X"00000000",
		16#6c85# => X"0001b20c",
		16#6c86# => X"0001b20c",
		16#6c87# => X"0001b214",
		16#6c88# => X"0001b214",
		16#6c89# => X"0001b21c",
		16#6c8a# => X"0001b21c",
		16#6c8b# => X"0001b224",
		16#6c8c# => X"0001b224",
		16#6c8d# => X"0001b22c",
		16#6c8e# => X"0001b22c",
		16#6c8f# => X"0001b234",
		16#6c90# => X"0001b234",
		16#6c91# => X"0001b23c",
		16#6c92# => X"0001b23c",
		16#6c93# => X"0001b244",
		16#6c94# => X"0001b244",
		16#6c95# => X"0001b24c",
		16#6c96# => X"0001b24c",
		16#6c97# => X"0001b254",
		16#6c98# => X"0001b254",
		16#6c99# => X"0001b25c",
		16#6c9a# => X"0001b25c",
		16#6c9b# => X"0001b264",
		16#6c9c# => X"0001b264",
		16#6c9d# => X"0001b26c",
		16#6c9e# => X"0001b26c",
		16#6c9f# => X"0001b274",
		16#6ca0# => X"0001b274",
		16#6ca1# => X"0001b27c",
		16#6ca2# => X"0001b27c",
		16#6ca3# => X"0001b284",
		16#6ca4# => X"0001b284",
		16#6ca5# => X"0001b28c",
		16#6ca6# => X"0001b28c",
		16#6ca7# => X"0001b294",
		16#6ca8# => X"0001b294",
		16#6ca9# => X"0001b29c",
		16#6caa# => X"0001b29c",
		16#6cab# => X"0001b2a4",
		16#6cac# => X"0001b2a4",
		16#6cad# => X"0001b2ac",
		16#6cae# => X"0001b2ac",
		16#6caf# => X"0001b2b4",
		16#6cb0# => X"0001b2b4",
		16#6cb1# => X"0001b2bc",
		16#6cb2# => X"0001b2bc",
		16#6cb3# => X"0001b2c4",
		16#6cb4# => X"0001b2c4",
		16#6cb5# => X"0001b2cc",
		16#6cb6# => X"0001b2cc",
		16#6cb7# => X"0001b2d4",
		16#6cb8# => X"0001b2d4",
		16#6cb9# => X"0001b2dc",
		16#6cba# => X"0001b2dc",
		16#6cbb# => X"0001b2e4",
		16#6cbc# => X"0001b2e4",
		16#6cbd# => X"0001b2ec",
		16#6cbe# => X"0001b2ec",
		16#6cbf# => X"0001b2f4",
		16#6cc0# => X"0001b2f4",
		16#6cc1# => X"0001b2fc",
		16#6cc2# => X"0001b2fc",
		16#6cc3# => X"0001b304",
		16#6cc4# => X"0001b304",
		16#6cc5# => X"0001b30c",
		16#6cc6# => X"0001b30c",
		16#6cc7# => X"0001b314",
		16#6cc8# => X"0001b314",
		16#6cc9# => X"0001b31c",
		16#6cca# => X"0001b31c",
		16#6ccb# => X"0001b324",
		16#6ccc# => X"0001b324",
		16#6ccd# => X"0001b32c",
		16#6cce# => X"0001b32c",
		16#6ccf# => X"0001b334",
		16#6cd0# => X"0001b334",
		16#6cd1# => X"0001b33c",
		16#6cd2# => X"0001b33c",
		16#6cd3# => X"0001b344",
		16#6cd4# => X"0001b344",
		16#6cd5# => X"0001b34c",
		16#6cd6# => X"0001b34c",
		16#6cd7# => X"0001b354",
		16#6cd8# => X"0001b354",
		16#6cd9# => X"0001b35c",
		16#6cda# => X"0001b35c",
		16#6cdb# => X"0001b364",
		16#6cdc# => X"0001b364",
		16#6cdd# => X"0001b36c",
		16#6cde# => X"0001b36c",
		16#6cdf# => X"0001b374",
		16#6ce0# => X"0001b374",
		16#6ce1# => X"0001b37c",
		16#6ce2# => X"0001b37c",
		16#6ce3# => X"0001b384",
		16#6ce4# => X"0001b384",
		16#6ce5# => X"0001b38c",
		16#6ce6# => X"0001b38c",
		16#6ce7# => X"0001b394",
		16#6ce8# => X"0001b394",
		16#6ce9# => X"0001b39c",
		16#6cea# => X"0001b39c",
		16#6ceb# => X"0001b3a4",
		16#6cec# => X"0001b3a4",
		16#6ced# => X"0001b3ac",
		16#6cee# => X"0001b3ac",
		16#6cef# => X"0001b3b4",
		16#6cf0# => X"0001b3b4",
		16#6cf1# => X"0001b3bc",
		16#6cf2# => X"0001b3bc",
		16#6cf3# => X"0001b3c4",
		16#6cf4# => X"0001b3c4",
		16#6cf5# => X"0001b3cc",
		16#6cf6# => X"0001b3cc",
		16#6cf7# => X"0001b3d4",
		16#6cf8# => X"0001b3d4",
		16#6cf9# => X"0001b3dc",
		16#6cfa# => X"0001b3dc",
		16#6cfb# => X"0001b3e4",
		16#6cfc# => X"0001b3e4",
		16#6cfd# => X"0001b3ec",
		16#6cfe# => X"0001b3ec",
		16#6cff# => X"0001b3f4",
		16#6d00# => X"0001b3f4",
		16#6d01# => X"0001b3fc",
		16#6d02# => X"0001b3fc",
		16#6d03# => X"0001b404",
		16#6d04# => X"0001b404",
		16#6d05# => X"0001b40c",
		16#6d06# => X"0001b40c",
		16#6d07# => X"0001b414",
		16#6d08# => X"0001b414",
		16#6d09# => X"0001b41c",
		16#6d0a# => X"0001b41c",
		16#6d0b# => X"0001b424",
		16#6d0c# => X"0001b424",
		16#6d0d# => X"0001b42c",
		16#6d0e# => X"0001b42c",
		16#6d0f# => X"0001b434",
		16#6d10# => X"0001b434",
		16#6d11# => X"0001b43c",
		16#6d12# => X"0001b43c",
		16#6d13# => X"0001b444",
		16#6d14# => X"0001b444",
		16#6d15# => X"0001b44c",
		16#6d16# => X"0001b44c",
		16#6d17# => X"0001b454",
		16#6d18# => X"0001b454",
		16#6d19# => X"0001b45c",
		16#6d1a# => X"0001b45c",
		16#6d1b# => X"0001b464",
		16#6d1c# => X"0001b464",
		16#6d1d# => X"0001b46c",
		16#6d1e# => X"0001b46c",
		16#6d1f# => X"0001b474",
		16#6d20# => X"0001b474",
		16#6d21# => X"0001b47c",
		16#6d22# => X"0001b47c",
		16#6d23# => X"0001b484",
		16#6d24# => X"0001b484",
		16#6d25# => X"0001b48c",
		16#6d26# => X"0001b48c",
		16#6d27# => X"0001b494",
		16#6d28# => X"0001b494",
		16#6d29# => X"0001b49c",
		16#6d2a# => X"0001b49c",
		16#6d2b# => X"0001b4a4",
		16#6d2c# => X"0001b4a4",
		16#6d2d# => X"0001b4ac",
		16#6d2e# => X"0001b4ac",
		16#6d2f# => X"0001b4b4",
		16#6d30# => X"0001b4b4",
		16#6d31# => X"0001b4bc",
		16#6d32# => X"0001b4bc",
		16#6d33# => X"0001b4c4",
		16#6d34# => X"0001b4c4",
		16#6d35# => X"0001b4cc",
		16#6d36# => X"0001b4cc",
		16#6d37# => X"0001b4d4",
		16#6d38# => X"0001b4d4",
		16#6d39# => X"0001b4dc",
		16#6d3a# => X"0001b4dc",
		16#6d3b# => X"0001b4e4",
		16#6d3c# => X"0001b4e4",
		16#6d3d# => X"0001b4ec",
		16#6d3e# => X"0001b4ec",
		16#6d3f# => X"0001b4f4",
		16#6d40# => X"0001b4f4",
		16#6d41# => X"0001b4fc",
		16#6d42# => X"0001b4fc",
		16#6d43# => X"0001b504",
		16#6d44# => X"0001b504",
		16#6d45# => X"0001b50c",
		16#6d46# => X"0001b50c",
		16#6d47# => X"0001b514",
		16#6d48# => X"0001b514",
		16#6d49# => X"0001b51c",
		16#6d4a# => X"0001b51c",
		16#6d4b# => X"0001b524",
		16#6d4c# => X"0001b524",
		16#6d4d# => X"0001b52c",
		16#6d4e# => X"0001b52c",
		16#6d4f# => X"0001b534",
		16#6d50# => X"0001b534",
		16#6d51# => X"0001b53c",
		16#6d52# => X"0001b53c",
		16#6d53# => X"0001b544",
		16#6d54# => X"0001b544",
		16#6d55# => X"0001b54c",
		16#6d56# => X"0001b54c",
		16#6d57# => X"0001b554",
		16#6d58# => X"0001b554",
		16#6d59# => X"0001b55c",
		16#6d5a# => X"0001b55c",
		16#6d5b# => X"0001b564",
		16#6d5c# => X"0001b564",
		16#6d5d# => X"0001b56c",
		16#6d5e# => X"0001b56c",
		16#6d5f# => X"0001b574",
		16#6d60# => X"0001b574",
		16#6d61# => X"0001b57c",
		16#6d62# => X"0001b57c",
		16#6d63# => X"0001b584",
		16#6d64# => X"0001b584",
		16#6d65# => X"0001b58c",
		16#6d66# => X"0001b58c",
		16#6d67# => X"0001b594",
		16#6d68# => X"0001b594",
		16#6d69# => X"0001b59c",
		16#6d6a# => X"0001b59c",
		16#6d6b# => X"0001b5a4",
		16#6d6c# => X"0001b5a4",
		16#6d6d# => X"0001b5ac",
		16#6d6e# => X"0001b5ac",
		16#6d6f# => X"0001b5b4",
		16#6d70# => X"0001b5b4",
		16#6d71# => X"0001b5bc",
		16#6d72# => X"0001b5bc",
		16#6d73# => X"0001b5c4",
		16#6d74# => X"0001b5c4",
		16#6d75# => X"0001b5cc",
		16#6d76# => X"0001b5cc",
		16#6d77# => X"0001b5d4",
		16#6d78# => X"0001b5d4",
		16#6d79# => X"0001b5dc",
		16#6d7a# => X"0001b5dc",
		16#6d7b# => X"0001b5e4",
		16#6d7c# => X"0001b5e4",
		16#6d7d# => X"0001b5ec",
		16#6d7e# => X"0001b5ec",
		16#6d7f# => X"0001b5f4",
		16#6d80# => X"0001b5f4",
		16#6d81# => X"0001b5fc",
		16#6d82# => X"0001b5fc",
		16#6d83# => X"0001b604",
		16#6d84# => X"0001b604",
		16#6d85# => X"00020000",
		16#6d86# => X"ffffffff",
		16#6d87# => X"ffffffff",
		16#6d88# => X"ffffffff",
		16#6d89# => X"ffffffff",
		16#6d8a# => X"ffffffff",
		16#6d8b# => X"ffffffff",
		16#6d8c# => X"ffffffff",
		16#6d8d# => X"ffffffff",
		16#6d8e# => X"ffffffff",
		16#6d8f# => X"ffffffff",
		16#6d90# => X"ffffffff",
		16#6d91# => X"ffffffff",
		16#6d92# => X"ffffffff",
		16#6d93# => X"ffffffff",
		16#6d94# => X"ffffffff",
		16#6d95# => X"ffffffff",
		16#6d96# => X"ffffffff",
		16#6d97# => X"ffffffff",
		16#6d98# => X"ffffffff",
		16#6d99# => X"ffffffff",
		16#6d9a# => X"ffffffff",
		16#6d9b# => X"ffffffff",
		16#6d9c# => X"ffffffff",
		16#6d9d# => X"ffffffff",
		16#6d9e# => X"ffffffff",
		16#6d9f# => X"ffffffff",
		16#6da0# => X"ffffffff",
		16#6da1# => X"ffffffff",
		16#6da2# => X"ffffffff",
		16#6da3# => X"ffffffff",
		16#6da4# => X"ffffffff",
		16#6da5# => X"ffffffff",
		16#6da6# => X"ffffffff",
		16#6da7# => X"ffffffff",
		16#6da8# => X"ffffffff",
		16#6da9# => X"ffffffff",
		16#6daa# => X"ffffffff",
		16#6dab# => X"ffffffff",
		16#6dac# => X"ffffffff",
		16#6dad# => X"ffffffff",
		16#6dae# => X"ffffffff",
		16#6daf# => X"ffffffff",
		16#6db0# => X"ffffffff",
		16#6db1# => X"ffffffff",
		16#6db2# => X"ffffffff",
		16#6db3# => X"ffffffff",
		16#6db4# => X"ffffffff",
		16#6db5# => X"ffffffff",
		16#6db6# => X"ffffffff",
		16#6db7# => X"ffffffff",
		16#6db8# => X"ffffffff",
		16#6db9# => X"ffffffff",
		16#6dba# => X"ffffffff",
		16#6dbb# => X"ffffffff",
		16#6dbc# => X"ffffffff",
		16#6dbd# => X"ffffffff",
		16#6dbe# => X"ffffffff",
		16#6dbf# => X"ffffffff",
		16#6dc0# => X"ffffffff",
		16#6dc1# => X"ffffffff",
		16#6dc2# => X"ffffffff",
		16#6dc3# => X"ffffffff",
		16#6dc4# => X"ffffffff",
		16#6dc5# => X"ffffffff",
		16#6dc6# => X"ffffffff",
		16#6dc7# => X"ffffffff",
		16#6dc8# => X"ffffffff",
		16#6dc9# => X"ffffffff",
		16#6dca# => X"ffffffff",
		16#6dcb# => X"ffffffff",
		16#6dcc# => X"ffffffff",
		16#6dcd# => X"ffffffff",
		16#6dce# => X"ffffffff",
		16#6dcf# => X"ffffffff",
		16#6dd0# => X"ffffffff",
		16#6dd1# => X"ffffffff",
		16#6dd2# => X"ffffffff",
		16#6dd3# => X"ffffffff",
		16#6dd4# => X"ffffffff",
		16#6dd5# => X"ffffffff",
		16#6dd6# => X"ffffffff",
		16#6dd7# => X"ffffffff",
		16#6dd8# => X"ffffffff",
		16#6dd9# => X"ffffffff",
		16#6dda# => X"ffffffff",
		16#6ddb# => X"ffffffff",
		16#6ddc# => X"ffffffff",
		16#6ddd# => X"ffffffff",
		16#6dde# => X"ffffffff",
		16#6ddf# => X"ffffffff",
		16#6de0# => X"ffffffff",
		16#6de1# => X"ffffffff",
		16#6de2# => X"ffffffff",
		16#6de3# => X"ffffffff",
		16#6de4# => X"00000001",
		16#6de5# => X"00000001",
		16#6de6# => X"41534349",
		16#6de7# => X"49000000",
		16#6de8# => X"00000000",
		16#6de9# => X"00000000",
		16#6dea# => X"00000000",
		16#6deb# => X"00000000",
		16#6dec# => X"00000000",
		16#6ded# => X"00000000",
		16#6dee# => X"41534349",
		16#6def# => X"49000000",
		16#6df0# => X"00000000",
		16#6df1# => X"00000000",
		16#6df2# => X"00000000",
		16#6df3# => X"00000000",
		16#6df4# => X"00000000",
		16#6df5# => X"00000000",
		16#6df6# => X"0001764c",
		16#6df7# => X"0001c50c",
		16#6df8# => X"00000000",
		others => X"00000000"
	);

end package;