library ieee;
use ieee.std_logic_1164.all;

package counter_config is

    constant CFG_COUNTER_N_COUNTER : integer range 1 to 16 := 4;

end package;

